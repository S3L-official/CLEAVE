module Cipher ( clk, rst, EncDec, Input, Key, Tweak, Output );
  input [63:0] Input;
  input [63:0] Key;
  output [63:0] Output;
  (* FIRMER="clock" *)input clk;
  (* FIRMER="control" *)input rst;
  (* FIRMER="control" *)input EncDec;
  wire   \MCInst_XOR_r0_Inst_0_n3 , \MCInst_XOR_r0_Inst_1_n3 ,
         \MCInst_XOR_r0_Inst_2_n3 , \MCInst_XOR_r0_Inst_3_n3 ,
         \MCInst_XOR_r0_Inst_4_n3 , \MCInst_XOR_r0_Inst_5_n3 ,
         \MCInst_XOR_r0_Inst_6_n3 , \MCInst_XOR_r0_Inst_7_n3 ,
         \MCInst_XOR_r0_Inst_8_n3 , \MCInst_XOR_r0_Inst_9_n3 ,
         \MCInst_XOR_r0_Inst_10_n3 , \MCInst_XOR_r0_Inst_11_n3 ,
         \MCInst_XOR_r0_Inst_12_n3 , \MCInst_XOR_r0_Inst_13_n3 ,
         \MCInst_XOR_r0_Inst_14_n3 , \MCInst_XOR_r0_Inst_15_n3 ,
         \AddKeyXOR1_XORInst_0_0_n2 , \AddKeyXOR1_XORInst_0_2_n2 ,
         \AddKeyXOR1_XORInst_1_0_n2 , \AddKeyXOR1_XORInst_1_2_n2 ,
         \AddKeyXOR1_XORInst_2_0_n2 , \AddKeyXOR1_XORInst_2_2_n2 ,
         \AddKeyXOR1_XORInst_3_0_n2 , \AddKeyXOR1_XORInst_3_2_n2 ,
         \AddKeyConstXOR_XORInst_0_0_n3 , \AddKeyConstXOR_XORInst_0_2_n3 ,
         \AddKeyConstXOR_XORInst_1_0_n3 , \AddKeyConstXOR_XORInst_1_2_n3 ,
         \AddKeyXOR2_XORInst_0_0_n2 , \AddKeyXOR2_XORInst_0_2_n2 ,
         \AddKeyXOR2_XORInst_1_0_n2 , \AddKeyXOR2_XORInst_1_2_n2 ,
         \AddKeyXOR2_XORInst_2_0_n2 , \AddKeyXOR2_XORInst_2_2_n2 ,
         \AddKeyXOR2_XORInst_3_0_n2 , \AddKeyXOR2_XORInst_3_2_n2 ,
         \AddKeyXOR2_XORInst_4_0_n2 , \AddKeyXOR2_XORInst_4_2_n2 ,
         \AddKeyXOR2_XORInst_5_0_n2 , \AddKeyXOR2_XORInst_5_2_n2 ,
         \AddKeyXOR2_XORInst_6_0_n2 , \AddKeyXOR2_XORInst_6_2_n2 ,
         \AddKeyXOR2_XORInst_7_0_n2 , \AddKeyXOR2_XORInst_7_2_n2 ,
         \AddKeyXOR2_XORInst_8_0_n2 , \AddKeyXOR2_XORInst_8_2_n2 ,
         \AddKeyXOR2_XORInst_9_0_n2 , \AddKeyXOR2_XORInst_9_2_n2 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n17 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n16 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n15 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n14 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n48 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n47 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n46 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n45 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n17 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n16 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n15 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n14 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n48 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n47 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n46 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n45 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n17 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n16 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n15 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n14 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n48 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n47 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n46 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n45 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n17 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n16 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n15 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n14 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n48 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n47 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n46 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n45 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n17 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n16 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n15 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n14 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n48 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n47 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n46 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n45 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n17 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n16 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n15 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n14 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n48 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n47 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n46 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n45 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n17 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n16 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n15 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n14 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n48 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n47 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n46 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n45 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n17 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n16 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n15 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n14 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n48 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n47 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n46 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n45 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n17 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n16 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n15 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n14 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n48 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n47 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n46 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n45 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n17 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n16 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n15 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n14 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n48 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n47 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n46 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n45 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n17 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n16 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n15 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n14 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n48 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n47 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n46 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n45 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n17 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n16 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n15 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n14 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n48 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n47 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n46 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n45 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n17 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n16 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n15 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n14 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n48 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n47 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n46 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n45 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n17 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n16 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n15 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n14 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n48 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n47 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n46 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n45 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n17 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n16 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n15 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n14 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n48 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n47 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n46 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n45 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n17 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n16 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n15 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n14 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n26 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n25 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n24 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n23 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n22 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n21 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n20 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n19 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n18 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n48 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n47 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n46 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n45 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n44 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n43 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n42 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n41 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n40 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n39 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n38 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n37 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n36 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n35 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n34 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n33 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n32 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n31 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n30 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n29 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n28 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n27 ,
         \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n26 ,
         \Red_PlaintextInst_LFInst_0_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_0_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_0_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_1_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_1_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_1_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_2_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_2_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_2_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_3_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_3_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_3_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_4_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_4_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_4_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_5_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_5_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_5_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_6_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_6_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_6_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_7_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_7_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_7_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_8_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_8_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_8_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_9_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_9_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_9_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_10_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_10_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_10_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_11_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_11_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_11_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_12_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_12_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_12_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_13_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_13_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_13_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_14_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_14_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_14_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_15_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_15_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_15_LFInst_2_n2 ,
         \Red_MCInst_XOR_r0_Inst_0_n3 , \Red_MCInst_XOR_r0_Inst_1_n3 ,
         \Red_MCInst_XOR_r0_Inst_2_n3 , \Red_MCInst_XOR_r0_Inst_3_n3 ,
         \Red_MCInst_XOR_r0_Inst_4_n3 , \Red_MCInst_XOR_r0_Inst_5_n3 ,
         \Red_MCInst_XOR_r0_Inst_6_n3 , \Red_MCInst_XOR_r0_Inst_7_n3 ,
         \Red_MCInst_XOR_r0_Inst_8_n3 , \Red_MCInst_XOR_r0_Inst_9_n3 ,
         \Red_MCInst_XOR_r0_Inst_10_n3 , \Red_MCInst_XOR_r0_Inst_11_n3 ,
         \StateRegOutputF_inst_LFInst_0_LFInst_0_n2 ,
         \StateRegOutputF_inst_LFInst_0_LFInst_1_n2 ,
         \StateRegOutputF_inst_LFInst_0_LFInst_2_n2 ,
         \StateRegOutputF_inst_LFInst_1_LFInst_0_n2 ,
         \StateRegOutputF_inst_LFInst_1_LFInst_1_n2 ,
         \StateRegOutputF_inst_LFInst_1_LFInst_2_n2 ,
         \StateRegOutputF_inst_LFInst_2_LFInst_0_n2 ,
         \StateRegOutputF_inst_LFInst_2_LFInst_1_n2 ,
         \StateRegOutputF_inst_LFInst_2_LFInst_2_n2 ,
         \StateRegOutputF_inst_LFInst_3_LFInst_0_n2 ,
         \StateRegOutputF_inst_LFInst_3_LFInst_1_n2 ,
         \StateRegOutputF_inst_LFInst_3_LFInst_2_n2 ,
         \StateRegOutputF_inst_LFInst_4_LFInst_0_n2 ,
         \StateRegOutputF_inst_LFInst_4_LFInst_1_n2 ,
         \StateRegOutputF_inst_LFInst_4_LFInst_2_n2 ,
         \StateRegOutputF_inst_LFInst_5_LFInst_0_n2 ,
         \StateRegOutputF_inst_LFInst_5_LFInst_1_n2 ,
         \StateRegOutputF_inst_LFInst_5_LFInst_2_n2 ,
         \StateRegOutputF_inst_LFInst_6_LFInst_0_n2 ,
         \StateRegOutputF_inst_LFInst_6_LFInst_1_n2 ,
         \StateRegOutputF_inst_LFInst_6_LFInst_2_n2 ,
         \StateRegOutputF_inst_LFInst_7_LFInst_0_n2 ,
         \StateRegOutputF_inst_LFInst_7_LFInst_1_n2 ,
         \StateRegOutputF_inst_LFInst_7_LFInst_2_n2 ,
         \StateRegOutputF_inst_LFInst_8_LFInst_0_n2 ,
         \StateRegOutputF_inst_LFInst_8_LFInst_1_n2 ,
         \StateRegOutputF_inst_LFInst_8_LFInst_2_n2 ,
         \StateRegOutputF_inst_LFInst_9_LFInst_0_n2 ,
         \StateRegOutputF_inst_LFInst_9_LFInst_1_n2 ,
         \StateRegOutputF_inst_LFInst_9_LFInst_2_n2 ,
         \StateRegOutputF_inst_LFInst_10_LFInst_0_n2 ,
         \StateRegOutputF_inst_LFInst_10_LFInst_1_n2 ,
         \StateRegOutputF_inst_LFInst_10_LFInst_2_n2 ,
         \StateRegOutputF_inst_LFInst_11_LFInst_0_n2 ,
         \StateRegOutputF_inst_LFInst_11_LFInst_1_n2 ,
         \StateRegOutputF_inst_LFInst_11_LFInst_2_n2 ,
         \StateRegOutputF_inst_LFInst_12_LFInst_0_n2 ,
         \StateRegOutputF_inst_LFInst_12_LFInst_1_n2 ,
         \StateRegOutputF_inst_LFInst_12_LFInst_2_n2 ,
         \StateRegOutputF_inst_LFInst_13_LFInst_0_n2 ,
         \StateRegOutputF_inst_LFInst_13_LFInst_1_n2 ,
         \StateRegOutputF_inst_LFInst_13_LFInst_2_n2 ,
         \StateRegOutputF_inst_LFInst_14_LFInst_0_n2 ,
         \StateRegOutputF_inst_LFInst_14_LFInst_1_n2 ,
         \StateRegOutputF_inst_LFInst_14_LFInst_2_n2 ,
         \StateRegOutputF_inst_LFInst_15_LFInst_0_n2 ,
         \StateRegOutputF_inst_LFInst_15_LFInst_1_n2 ,
         \StateRegOutputF_inst_LFInst_15_LFInst_2_n2 ,
         \CipherErrorVecGen_XORInst_0_0_n4 ,
         \CipherErrorVecGen_XORInst_0_1_n2 ,
         \CipherErrorVecGen_XORInst_0_2_n3 ,
         \CipherErrorVecGen_XORInst_1_0_n4 ,
         \CipherErrorVecGen_XORInst_1_1_n2 ,
         \CipherErrorVecGen_XORInst_1_2_n3 ,
         \CipherErrorVecGen_XORInst_2_0_n4 ,
         \CipherErrorVecGen_XORInst_2_1_n2 ,
         \CipherErrorVecGen_XORInst_2_2_n3 ,
         \CipherErrorVecGen_XORInst_3_0_n4 ,
         \CipherErrorVecGen_XORInst_3_1_n2 ,
         \CipherErrorVecGen_XORInst_3_2_n3 ,
         \CipherErrorVecGen_XORInst_4_0_n4 ,
         \CipherErrorVecGen_XORInst_4_1_n2 ,
         \CipherErrorVecGen_XORInst_4_2_n3 ,
         \CipherErrorVecGen_XORInst_5_0_n4 ,
         \CipherErrorVecGen_XORInst_5_1_n2 ,
         \CipherErrorVecGen_XORInst_5_2_n3 ,
         \CipherErrorVecGen_XORInst_6_0_n4 ,
         \CipherErrorVecGen_XORInst_6_1_n2 ,
         \CipherErrorVecGen_XORInst_6_2_n3 ,
         \CipherErrorVecGen_XORInst_7_0_n4 ,
         \CipherErrorVecGen_XORInst_7_1_n2 ,
         \CipherErrorVecGen_XORInst_7_2_n3 ,
         \CipherErrorVecGen_XORInst_8_0_n4 ,
         \CipherErrorVecGen_XORInst_8_1_n2 ,
         \CipherErrorVecGen_XORInst_8_2_n3 ,
         \CipherErrorVecGen_XORInst_9_0_n4 ,
         \CipherErrorVecGen_XORInst_9_1_n2 ,
         \CipherErrorVecGen_XORInst_9_2_n3 ,
         \CipherErrorVecGen_XORInst_10_0_n4 ,
         \CipherErrorVecGen_XORInst_10_1_n2 ,
         \CipherErrorVecGen_XORInst_10_2_n3 ,
         \CipherErrorVecGen_XORInst_11_0_n4 ,
         \CipherErrorVecGen_XORInst_11_1_n2 ,
         \CipherErrorVecGen_XORInst_11_2_n3 ,
         \CipherErrorVecGen_XORInst_12_0_n4 ,
         \CipherErrorVecGen_XORInst_12_1_n2 ,
         \CipherErrorVecGen_XORInst_12_2_n3 ,
         \CipherErrorVecGen_XORInst_13_0_n4 ,
         \CipherErrorVecGen_XORInst_13_1_n2 ,
         \CipherErrorVecGen_XORInst_13_2_n3 ,
         \CipherErrorVecGen_XORInst_14_0_n4 ,
         \CipherErrorVecGen_XORInst_14_1_n2 ,
         \CipherErrorVecGen_XORInst_14_2_n3 ,
         \CipherErrorVecGen_XORInst_15_0_n4 ,
         \CipherErrorVecGen_XORInst_15_1_n2 ,
         \CipherErrorVecGen_XORInst_15_2_n3 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n19 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n19 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n19 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n19 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n19 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n19 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n19 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n19 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n19 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n19 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n19 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n19 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n19 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n19 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n19 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n20 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n19 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n37 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n36 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n35 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n34 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n33 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n32 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n31 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n30 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n29 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n28 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n27 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n26 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n25 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n24 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n23 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n22 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n21 ,
         \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n20 ,
         \StateRegOutputF_inst2_LFInst_0_LFInst_0_n2 ,
         \StateRegOutputF_inst2_LFInst_0_LFInst_1_n2 ,
         \StateRegOutputF_inst2_LFInst_0_LFInst_2_n2 ,
         \StateRegOutputF_inst2_LFInst_1_LFInst_0_n2 ,
         \StateRegOutputF_inst2_LFInst_1_LFInst_1_n2 ,
         \StateRegOutputF_inst2_LFInst_1_LFInst_2_n2 ,
         \StateRegOutputF_inst2_LFInst_2_LFInst_0_n2 ,
         \StateRegOutputF_inst2_LFInst_2_LFInst_1_n2 ,
         \StateRegOutputF_inst2_LFInst_2_LFInst_2_n2 ,
         \StateRegOutputF_inst2_LFInst_3_LFInst_0_n2 ,
         \StateRegOutputF_inst2_LFInst_3_LFInst_1_n2 ,
         \StateRegOutputF_inst2_LFInst_3_LFInst_2_n2 ,
         \StateRegOutputF_inst2_LFInst_4_LFInst_0_n2 ,
         \StateRegOutputF_inst2_LFInst_4_LFInst_1_n2 ,
         \StateRegOutputF_inst2_LFInst_4_LFInst_2_n2 ,
         \StateRegOutputF_inst2_LFInst_5_LFInst_0_n2 ,
         \StateRegOutputF_inst2_LFInst_5_LFInst_1_n2 ,
         \StateRegOutputF_inst2_LFInst_5_LFInst_2_n2 ,
         \StateRegOutputF_inst2_LFInst_6_LFInst_0_n2 ,
         \StateRegOutputF_inst2_LFInst_6_LFInst_1_n2 ,
         \StateRegOutputF_inst2_LFInst_6_LFInst_2_n2 ,
         \StateRegOutputF_inst2_LFInst_7_LFInst_0_n2 ,
         \StateRegOutputF_inst2_LFInst_7_LFInst_1_n2 ,
         \StateRegOutputF_inst2_LFInst_7_LFInst_2_n2 ,
         \StateRegOutputF_inst2_LFInst_8_LFInst_0_n2 ,
         \StateRegOutputF_inst2_LFInst_8_LFInst_1_n2 ,
         \StateRegOutputF_inst2_LFInst_8_LFInst_2_n2 ,
         \StateRegOutputF_inst2_LFInst_9_LFInst_0_n2 ,
         \StateRegOutputF_inst2_LFInst_9_LFInst_1_n2 ,
         \StateRegOutputF_inst2_LFInst_9_LFInst_2_n2 ,
         \StateRegOutputF_inst2_LFInst_10_LFInst_0_n2 ,
         \StateRegOutputF_inst2_LFInst_10_LFInst_1_n2 ,
         \StateRegOutputF_inst2_LFInst_10_LFInst_2_n2 ,
         \StateRegOutputF_inst2_LFInst_11_LFInst_0_n2 ,
         \StateRegOutputF_inst2_LFInst_11_LFInst_1_n2 ,
         \StateRegOutputF_inst2_LFInst_11_LFInst_2_n2 ,
         \StateRegOutputF_inst2_LFInst_12_LFInst_0_n2 ,
         \StateRegOutputF_inst2_LFInst_12_LFInst_1_n2 ,
         \StateRegOutputF_inst2_LFInst_12_LFInst_2_n2 ,
         \StateRegOutputF_inst2_LFInst_13_LFInst_0_n2 ,
         \StateRegOutputF_inst2_LFInst_13_LFInst_1_n2 ,
         \StateRegOutputF_inst2_LFInst_13_LFInst_2_n2 ,
         \StateRegOutputF_inst2_LFInst_14_LFInst_0_n2 ,
         \StateRegOutputF_inst2_LFInst_14_LFInst_1_n2 ,
         \StateRegOutputF_inst2_LFInst_14_LFInst_2_n2 ,
         \StateRegOutputF_inst2_LFInst_15_LFInst_0_n2 ,
         \StateRegOutputF_inst2_LFInst_15_LFInst_1_n2 ,
         \StateRegOutputF_inst2_LFInst_15_LFInst_2_n2 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n27 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n26 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n25 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n24 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n23 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n22 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n21 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n20 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n27 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n26 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n25 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n24 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n23 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n22 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n21 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n20 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n27 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n26 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n25 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n24 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n23 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n22 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n21 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n20 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n27 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n26 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n25 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n24 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n23 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n22 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n21 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n20 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n27 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n26 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n25 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n24 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n23 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n22 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n21 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n20 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n27 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n26 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n25 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n24 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n23 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n22 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n21 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n20 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n27 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n26 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n25 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n24 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n23 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n22 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n21 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n20 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n27 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n26 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n25 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n24 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n23 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n22 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n21 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n20 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n27 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n26 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n25 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n24 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n23 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n22 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n21 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n20 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n27 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n26 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n25 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n24 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n23 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n22 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n21 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n20 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n27 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n26 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n25 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n24 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n23 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n22 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n21 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n20 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n27 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n26 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n25 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n24 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n23 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n22 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n21 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n20 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n27 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n26 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n25 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n24 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n23 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n22 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n21 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n20 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n27 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n26 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n25 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n24 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n23 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n22 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n21 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n20 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n27 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n26 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n25 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n24 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n23 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n22 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n21 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n20 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n27 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n26 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n25 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n24 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n23 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n22 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n21 ,
         \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n20 ,
         \Red_K0Inst_LFInst_0_LFInst_0_n2 , \Red_K0Inst_LFInst_0_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_0_LFInst_2_n2 , \Red_K0Inst_LFInst_1_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_1_LFInst_1_n2 , \Red_K0Inst_LFInst_1_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_2_LFInst_0_n2 , \Red_K0Inst_LFInst_2_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_2_LFInst_2_n2 , \Red_K0Inst_LFInst_3_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_3_LFInst_1_n2 , \Red_K0Inst_LFInst_3_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_4_LFInst_0_n2 , \Red_K0Inst_LFInst_4_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_4_LFInst_2_n2 , \Red_K0Inst_LFInst_5_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_5_LFInst_1_n2 , \Red_K0Inst_LFInst_5_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_6_LFInst_0_n2 , \Red_K0Inst_LFInst_6_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_6_LFInst_2_n2 , \Red_K0Inst_LFInst_7_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_7_LFInst_1_n2 , \Red_K0Inst_LFInst_7_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_8_LFInst_0_n2 , \Red_K0Inst_LFInst_8_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_8_LFInst_2_n2 , \Red_K0Inst_LFInst_9_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_9_LFInst_1_n2 , \Red_K0Inst_LFInst_9_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_10_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_10_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_10_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_11_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_11_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_11_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_12_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_12_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_12_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_13_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_13_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_13_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_14_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_14_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_14_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_15_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_15_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_15_LFInst_2_n2 ;
  wire   [63:0] MCOutput;
  wire   [63:0] AddRoundKeyOutput;
  wire   [47:0] CipherErrorVec;
  wire   [63:0] PermutationInput;
  wire   [63:0] Feedback;
  wire   [47:0] Red_Input;
  wire   [47:0] Red_MCOutput;
  wire   [47:0] Red_K0;
  wire   [47:0] Red_AddRoundKeyOutput;
  wire   [47:0] StateRegOutputF;
  wire   [47:0] Red_PermutationInput;
  wire   [47:0] Red_Feedback;
  wire   [47:0] FeedbackF;
  wire   [47:0] CipherErrorVec2;

  XNOR2_X1 \MCInst_XOR_r0_Inst_0_U2  ( .A(\MCInst_XOR_r0_Inst_0_n3 ), .B(
        Input[0]), .ZN(MCOutput[48]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_0_U1  ( .A(Input[48]), .B(Input[16]), .ZN(
        \MCInst_XOR_r0_Inst_0_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_0_U1  ( .A(Input[32]), .B(Input[0]), .Z(
        MCOutput[32]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_1_U2  ( .A(\MCInst_XOR_r0_Inst_1_n3 ), .B(
        Input[1]), .ZN(MCOutput[49]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_1_U1  ( .A(Input[49]), .B(Input[17]), .ZN(
        \MCInst_XOR_r0_Inst_1_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_1_U1  ( .A(Input[33]), .B(Input[1]), .Z(
        MCOutput[33]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_2_U2  ( .A(\MCInst_XOR_r0_Inst_2_n3 ), .B(
        Input[2]), .ZN(MCOutput[50]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_2_U1  ( .A(Input[50]), .B(Input[18]), .ZN(
        \MCInst_XOR_r0_Inst_2_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_2_U1  ( .A(Input[34]), .B(Input[2]), .Z(
        MCOutput[34]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_3_U2  ( .A(\MCInst_XOR_r0_Inst_3_n3 ), .B(
        Input[3]), .ZN(MCOutput[51]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_3_U1  ( .A(Input[51]), .B(Input[19]), .ZN(
        \MCInst_XOR_r0_Inst_3_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_3_U1  ( .A(Input[35]), .B(Input[3]), .Z(
        MCOutput[35]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_4_U2  ( .A(\MCInst_XOR_r0_Inst_4_n3 ), .B(
        Input[4]), .ZN(MCOutput[52]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_4_U1  ( .A(Input[52]), .B(Input[20]), .ZN(
        \MCInst_XOR_r0_Inst_4_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_4_U1  ( .A(Input[36]), .B(Input[4]), .Z(
        MCOutput[36]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_5_U2  ( .A(\MCInst_XOR_r0_Inst_5_n3 ), .B(
        Input[5]), .ZN(MCOutput[53]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_5_U1  ( .A(Input[53]), .B(Input[21]), .ZN(
        \MCInst_XOR_r0_Inst_5_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_5_U1  ( .A(Input[37]), .B(Input[5]), .Z(
        MCOutput[37]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_6_U2  ( .A(\MCInst_XOR_r0_Inst_6_n3 ), .B(
        Input[6]), .ZN(MCOutput[54]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_6_U1  ( .A(Input[54]), .B(Input[22]), .ZN(
        \MCInst_XOR_r0_Inst_6_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_6_U1  ( .A(Input[38]), .B(Input[6]), .Z(
        MCOutput[38]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_7_U2  ( .A(\MCInst_XOR_r0_Inst_7_n3 ), .B(
        Input[7]), .ZN(MCOutput[55]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_7_U1  ( .A(Input[55]), .B(Input[23]), .ZN(
        \MCInst_XOR_r0_Inst_7_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_7_U1  ( .A(Input[39]), .B(Input[7]), .Z(
        MCOutput[39]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_8_U2  ( .A(\MCInst_XOR_r0_Inst_8_n3 ), .B(
        Input[8]), .ZN(MCOutput[56]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_8_U1  ( .A(Input[56]), .B(Input[24]), .ZN(
        \MCInst_XOR_r0_Inst_8_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_8_U1  ( .A(Input[40]), .B(Input[8]), .Z(
        MCOutput[40]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_9_U2  ( .A(\MCInst_XOR_r0_Inst_9_n3 ), .B(
        Input[9]), .ZN(MCOutput[57]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_9_U1  ( .A(Input[57]), .B(Input[25]), .ZN(
        \MCInst_XOR_r0_Inst_9_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_9_U1  ( .A(Input[41]), .B(Input[9]), .Z(
        MCOutput[41]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_10_U2  ( .A(\MCInst_XOR_r0_Inst_10_n3 ), .B(
        Input[10]), .ZN(MCOutput[58]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_10_U1  ( .A(Input[58]), .B(Input[26]), .ZN(
        \MCInst_XOR_r0_Inst_10_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_10_U1  ( .A(Input[42]), .B(Input[10]), .Z(
        MCOutput[42]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_11_U2  ( .A(\MCInst_XOR_r0_Inst_11_n3 ), .B(
        Input[11]), .ZN(MCOutput[59]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_11_U1  ( .A(Input[59]), .B(Input[27]), .ZN(
        \MCInst_XOR_r0_Inst_11_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_11_U1  ( .A(Input[43]), .B(Input[11]), .Z(
        MCOutput[43]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_12_U2  ( .A(\MCInst_XOR_r0_Inst_12_n3 ), .B(
        Input[12]), .ZN(MCOutput[60]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_12_U1  ( .A(Input[60]), .B(Input[28]), .ZN(
        \MCInst_XOR_r0_Inst_12_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_12_U1  ( .A(Input[44]), .B(Input[12]), .Z(
        MCOutput[44]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_13_U2  ( .A(\MCInst_XOR_r0_Inst_13_n3 ), .B(
        Input[13]), .ZN(MCOutput[61]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_13_U1  ( .A(Input[61]), .B(Input[29]), .ZN(
        \MCInst_XOR_r0_Inst_13_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_13_U1  ( .A(Input[45]), .B(Input[13]), .Z(
        MCOutput[45]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_14_U2  ( .A(\MCInst_XOR_r0_Inst_14_n3 ), .B(
        Input[14]), .ZN(MCOutput[62]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_14_U1  ( .A(Input[62]), .B(Input[30]), .ZN(
        \MCInst_XOR_r0_Inst_14_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_14_U1  ( .A(Input[46]), .B(Input[14]), .Z(
        MCOutput[46]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_15_U2  ( .A(\MCInst_XOR_r0_Inst_15_n3 ), .B(
        Input[15]), .ZN(MCOutput[63]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_15_U1  ( .A(Input[63]), .B(Input[31]), .ZN(
        \MCInst_XOR_r0_Inst_15_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_15_U1  ( .A(Input[47]), .B(Input[15]), .Z(
        MCOutput[47]) );
  INV_X1 \AddKeyXOR1_XORInst_0_0_U2  ( .A(\AddKeyXOR1_XORInst_0_0_n2 ), .ZN(
        AddRoundKeyOutput[48]) );
  XNOR2_X1 \AddKeyXOR1_XORInst_0_0_U1  ( .A(MCOutput[48]), .B(Key[48]), .ZN(
        \AddKeyXOR1_XORInst_0_0_n2 ) );
  XOR2_X2 \AddKeyXOR1_XORInst_0_1_U1  ( .A(MCOutput[49]), .B(Key[49]), .Z(
        AddRoundKeyOutput[49]) );
  INV_X1 \AddKeyXOR1_XORInst_0_2_U2  ( .A(\AddKeyXOR1_XORInst_0_2_n2 ), .ZN(
        AddRoundKeyOutput[50]) );
  XNOR2_X1 \AddKeyXOR1_XORInst_0_2_U1  ( .A(MCOutput[50]), .B(Key[50]), .ZN(
        \AddKeyXOR1_XORInst_0_2_n2 ) );
  XOR2_X2 \AddKeyXOR1_XORInst_0_3_U1  ( .A(MCOutput[51]), .B(Key[51]), .Z(
        AddRoundKeyOutput[51]) );
  INV_X1 \AddKeyXOR1_XORInst_1_0_U2  ( .A(\AddKeyXOR1_XORInst_1_0_n2 ), .ZN(
        AddRoundKeyOutput[52]) );
  XNOR2_X1 \AddKeyXOR1_XORInst_1_0_U1  ( .A(MCOutput[52]), .B(Key[52]), .ZN(
        \AddKeyXOR1_XORInst_1_0_n2 ) );
  XOR2_X2 \AddKeyXOR1_XORInst_1_1_U1  ( .A(MCOutput[53]), .B(Key[53]), .Z(
        AddRoundKeyOutput[53]) );
  INV_X1 \AddKeyXOR1_XORInst_1_2_U2  ( .A(\AddKeyXOR1_XORInst_1_2_n2 ), .ZN(
        AddRoundKeyOutput[54]) );
  XNOR2_X1 \AddKeyXOR1_XORInst_1_2_U1  ( .A(MCOutput[54]), .B(Key[54]), .ZN(
        \AddKeyXOR1_XORInst_1_2_n2 ) );
  XOR2_X2 \AddKeyXOR1_XORInst_1_3_U1  ( .A(MCOutput[55]), .B(Key[55]), .Z(
        AddRoundKeyOutput[55]) );
  INV_X1 \AddKeyXOR1_XORInst_2_0_U2  ( .A(\AddKeyXOR1_XORInst_2_0_n2 ), .ZN(
        AddRoundKeyOutput[56]) );
  XNOR2_X1 \AddKeyXOR1_XORInst_2_0_U1  ( .A(MCOutput[56]), .B(Key[56]), .ZN(
        \AddKeyXOR1_XORInst_2_0_n2 ) );
  XOR2_X2 \AddKeyXOR1_XORInst_2_1_U1  ( .A(MCOutput[57]), .B(Key[57]), .Z(
        AddRoundKeyOutput[57]) );
  INV_X1 \AddKeyXOR1_XORInst_2_2_U2  ( .A(\AddKeyXOR1_XORInst_2_2_n2 ), .ZN(
        AddRoundKeyOutput[58]) );
  XNOR2_X1 \AddKeyXOR1_XORInst_2_2_U1  ( .A(MCOutput[58]), .B(Key[58]), .ZN(
        \AddKeyXOR1_XORInst_2_2_n2 ) );
  XOR2_X2 \AddKeyXOR1_XORInst_2_3_U1  ( .A(MCOutput[59]), .B(Key[59]), .Z(
        AddRoundKeyOutput[59]) );
  INV_X1 \AddKeyXOR1_XORInst_3_0_U2  ( .A(\AddKeyXOR1_XORInst_3_0_n2 ), .ZN(
        AddRoundKeyOutput[60]) );
  XNOR2_X1 \AddKeyXOR1_XORInst_3_0_U1  ( .A(MCOutput[60]), .B(Key[60]), .ZN(
        \AddKeyXOR1_XORInst_3_0_n2 ) );
  XOR2_X2 \AddKeyXOR1_XORInst_3_1_U1  ( .A(MCOutput[61]), .B(Key[61]), .Z(
        AddRoundKeyOutput[61]) );
  INV_X1 \AddKeyXOR1_XORInst_3_2_U2  ( .A(\AddKeyXOR1_XORInst_3_2_n2 ), .ZN(
        AddRoundKeyOutput[62]) );
  XNOR2_X1 \AddKeyXOR1_XORInst_3_2_U1  ( .A(MCOutput[62]), .B(Key[62]), .ZN(
        \AddKeyXOR1_XORInst_3_2_n2 ) );
  XOR2_X2 \AddKeyXOR1_XORInst_3_3_U1  ( .A(MCOutput[63]), .B(Key[63]), .Z(
        AddRoundKeyOutput[63]) );
  INV_X1 \AddKeyConstXOR_XORInst_0_0_U2  ( .A(\AddKeyConstXOR_XORInst_0_0_n3 ), 
        .ZN(AddRoundKeyOutput[40]) );
  XNOR2_X1 \AddKeyConstXOR_XORInst_0_0_U1  ( .A(Key[40]), .B(MCOutput[40]), 
        .ZN(\AddKeyConstXOR_XORInst_0_0_n3 ) );
  XOR2_X2 \AddKeyConstXOR_XORInst_0_1_U1  ( .A(Key[41]), .B(MCOutput[41]), .Z(
        AddRoundKeyOutput[41]) );
  INV_X1 \AddKeyConstXOR_XORInst_0_2_U2  ( .A(\AddKeyConstXOR_XORInst_0_2_n3 ), 
        .ZN(AddRoundKeyOutput[42]) );
  XNOR2_X1 \AddKeyConstXOR_XORInst_0_2_U1  ( .A(Key[42]), .B(MCOutput[42]), 
        .ZN(\AddKeyConstXOR_XORInst_0_2_n3 ) );
  XOR2_X2 \AddKeyConstXOR_XORInst_0_3_U1  ( .A(Key[43]), .B(MCOutput[43]), .Z(
        AddRoundKeyOutput[43]) );
  INV_X1 \AddKeyConstXOR_XORInst_1_0_U2  ( .A(\AddKeyConstXOR_XORInst_1_0_n3 ), 
        .ZN(AddRoundKeyOutput[44]) );
  XNOR2_X1 \AddKeyConstXOR_XORInst_1_0_U1  ( .A(Key[44]), .B(MCOutput[44]), 
        .ZN(\AddKeyConstXOR_XORInst_1_0_n3 ) );
  XOR2_X2 \AddKeyConstXOR_XORInst_1_1_U1  ( .A(Key[45]), .B(MCOutput[45]), .Z(
        AddRoundKeyOutput[45]) );
  INV_X1 \AddKeyConstXOR_XORInst_1_2_U2  ( .A(\AddKeyConstXOR_XORInst_1_2_n3 ), 
        .ZN(AddRoundKeyOutput[46]) );
  XNOR2_X1 \AddKeyConstXOR_XORInst_1_2_U1  ( .A(Key[46]), .B(MCOutput[46]), 
        .ZN(\AddKeyConstXOR_XORInst_1_2_n3 ) );
  XOR2_X2 \AddKeyConstXOR_XORInst_1_3_U1  ( .A(Key[47]), .B(MCOutput[47]), .Z(
        AddRoundKeyOutput[47]) );
  INV_X1 \AddKeyXOR2_XORInst_0_0_U2  ( .A(\AddKeyXOR2_XORInst_0_0_n2 ), .ZN(
        AddRoundKeyOutput[0]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_0_0_U1  ( .A(Input[0]), .B(Key[0]), .ZN(
        \AddKeyXOR2_XORInst_0_0_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_0_1_U1  ( .A(Input[1]), .B(Key[1]), .Z(
        AddRoundKeyOutput[1]) );
  INV_X1 \AddKeyXOR2_XORInst_0_2_U2  ( .A(\AddKeyXOR2_XORInst_0_2_n2 ), .ZN(
        AddRoundKeyOutput[2]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_0_2_U1  ( .A(Input[2]), .B(Key[2]), .ZN(
        \AddKeyXOR2_XORInst_0_2_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_0_3_U1  ( .A(Input[3]), .B(Key[3]), .Z(
        AddRoundKeyOutput[3]) );
  INV_X1 \AddKeyXOR2_XORInst_1_0_U2  ( .A(\AddKeyXOR2_XORInst_1_0_n2 ), .ZN(
        AddRoundKeyOutput[4]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_1_0_U1  ( .A(Input[4]), .B(Key[4]), .ZN(
        \AddKeyXOR2_XORInst_1_0_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_1_1_U1  ( .A(Input[5]), .B(Key[5]), .Z(
        AddRoundKeyOutput[5]) );
  INV_X1 \AddKeyXOR2_XORInst_1_2_U2  ( .A(\AddKeyXOR2_XORInst_1_2_n2 ), .ZN(
        AddRoundKeyOutput[6]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_1_2_U1  ( .A(Input[6]), .B(Key[6]), .ZN(
        \AddKeyXOR2_XORInst_1_2_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_1_3_U1  ( .A(Input[7]), .B(Key[7]), .Z(
        AddRoundKeyOutput[7]) );
  INV_X1 \AddKeyXOR2_XORInst_2_0_U2  ( .A(\AddKeyXOR2_XORInst_2_0_n2 ), .ZN(
        AddRoundKeyOutput[8]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_2_0_U1  ( .A(Input[8]), .B(Key[8]), .ZN(
        \AddKeyXOR2_XORInst_2_0_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_2_1_U1  ( .A(Input[9]), .B(Key[9]), .Z(
        AddRoundKeyOutput[9]) );
  INV_X1 \AddKeyXOR2_XORInst_2_2_U2  ( .A(\AddKeyXOR2_XORInst_2_2_n2 ), .ZN(
        AddRoundKeyOutput[10]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_2_2_U1  ( .A(Input[10]), .B(Key[10]), .ZN(
        \AddKeyXOR2_XORInst_2_2_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_2_3_U1  ( .A(Input[11]), .B(Key[11]), .Z(
        AddRoundKeyOutput[11]) );
  INV_X1 \AddKeyXOR2_XORInst_3_0_U2  ( .A(\AddKeyXOR2_XORInst_3_0_n2 ), .ZN(
        AddRoundKeyOutput[12]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_3_0_U1  ( .A(Input[12]), .B(Key[12]), .ZN(
        \AddKeyXOR2_XORInst_3_0_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_3_1_U1  ( .A(Input[13]), .B(Key[13]), .Z(
        AddRoundKeyOutput[13]) );
  INV_X1 \AddKeyXOR2_XORInst_3_2_U2  ( .A(\AddKeyXOR2_XORInst_3_2_n2 ), .ZN(
        AddRoundKeyOutput[14]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_3_2_U1  ( .A(Input[14]), .B(Key[14]), .ZN(
        \AddKeyXOR2_XORInst_3_2_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_3_3_U1  ( .A(Input[15]), .B(Key[15]), .Z(
        AddRoundKeyOutput[15]) );
  INV_X1 \AddKeyXOR2_XORInst_4_0_U2  ( .A(\AddKeyXOR2_XORInst_4_0_n2 ), .ZN(
        AddRoundKeyOutput[16]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_4_0_U1  ( .A(Input[16]), .B(Key[16]), .ZN(
        \AddKeyXOR2_XORInst_4_0_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_4_1_U1  ( .A(Input[17]), .B(Key[17]), .Z(
        AddRoundKeyOutput[17]) );
  INV_X1 \AddKeyXOR2_XORInst_4_2_U2  ( .A(\AddKeyXOR2_XORInst_4_2_n2 ), .ZN(
        AddRoundKeyOutput[18]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_4_2_U1  ( .A(Input[18]), .B(Key[18]), .ZN(
        \AddKeyXOR2_XORInst_4_2_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_4_3_U1  ( .A(Input[19]), .B(Key[19]), .Z(
        AddRoundKeyOutput[19]) );
  INV_X1 \AddKeyXOR2_XORInst_5_0_U2  ( .A(\AddKeyXOR2_XORInst_5_0_n2 ), .ZN(
        AddRoundKeyOutput[20]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_5_0_U1  ( .A(Input[20]), .B(Key[20]), .ZN(
        \AddKeyXOR2_XORInst_5_0_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_5_1_U1  ( .A(Input[21]), .B(Key[21]), .Z(
        AddRoundKeyOutput[21]) );
  INV_X1 \AddKeyXOR2_XORInst_5_2_U2  ( .A(\AddKeyXOR2_XORInst_5_2_n2 ), .ZN(
        AddRoundKeyOutput[22]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_5_2_U1  ( .A(Input[22]), .B(Key[22]), .ZN(
        \AddKeyXOR2_XORInst_5_2_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_5_3_U1  ( .A(Input[23]), .B(Key[23]), .Z(
        AddRoundKeyOutput[23]) );
  INV_X1 \AddKeyXOR2_XORInst_6_0_U2  ( .A(\AddKeyXOR2_XORInst_6_0_n2 ), .ZN(
        AddRoundKeyOutput[24]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_6_0_U1  ( .A(Input[24]), .B(Key[24]), .ZN(
        \AddKeyXOR2_XORInst_6_0_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_6_1_U1  ( .A(Input[25]), .B(Key[25]), .Z(
        AddRoundKeyOutput[25]) );
  INV_X1 \AddKeyXOR2_XORInst_6_2_U2  ( .A(\AddKeyXOR2_XORInst_6_2_n2 ), .ZN(
        AddRoundKeyOutput[26]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_6_2_U1  ( .A(Input[26]), .B(Key[26]), .ZN(
        \AddKeyXOR2_XORInst_6_2_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_6_3_U1  ( .A(Input[27]), .B(Key[27]), .Z(
        AddRoundKeyOutput[27]) );
  INV_X1 \AddKeyXOR2_XORInst_7_0_U2  ( .A(\AddKeyXOR2_XORInst_7_0_n2 ), .ZN(
        AddRoundKeyOutput[28]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_7_0_U1  ( .A(Input[28]), .B(Key[28]), .ZN(
        \AddKeyXOR2_XORInst_7_0_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_7_1_U1  ( .A(Input[29]), .B(Key[29]), .Z(
        AddRoundKeyOutput[29]) );
  INV_X1 \AddKeyXOR2_XORInst_7_2_U2  ( .A(\AddKeyXOR2_XORInst_7_2_n2 ), .ZN(
        AddRoundKeyOutput[30]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_7_2_U1  ( .A(Input[30]), .B(Key[30]), .ZN(
        \AddKeyXOR2_XORInst_7_2_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_7_3_U1  ( .A(Input[31]), .B(Key[31]), .Z(
        AddRoundKeyOutput[31]) );
  INV_X1 \AddKeyXOR2_XORInst_8_0_U2  ( .A(\AddKeyXOR2_XORInst_8_0_n2 ), .ZN(
        AddRoundKeyOutput[32]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_8_0_U1  ( .A(MCOutput[32]), .B(Key[32]), .ZN(
        \AddKeyXOR2_XORInst_8_0_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_8_1_U1  ( .A(MCOutput[33]), .B(Key[33]), .Z(
        AddRoundKeyOutput[33]) );
  INV_X1 \AddKeyXOR2_XORInst_8_2_U2  ( .A(\AddKeyXOR2_XORInst_8_2_n2 ), .ZN(
        AddRoundKeyOutput[34]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_8_2_U1  ( .A(MCOutput[34]), .B(Key[34]), .ZN(
        \AddKeyXOR2_XORInst_8_2_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_8_3_U1  ( .A(MCOutput[35]), .B(Key[35]), .Z(
        AddRoundKeyOutput[35]) );
  INV_X1 \AddKeyXOR2_XORInst_9_0_U2  ( .A(\AddKeyXOR2_XORInst_9_0_n2 ), .ZN(
        AddRoundKeyOutput[36]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_9_0_U1  ( .A(MCOutput[36]), .B(Key[36]), .ZN(
        \AddKeyXOR2_XORInst_9_0_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_9_1_U1  ( .A(MCOutput[37]), .B(Key[37]), .Z(
        AddRoundKeyOutput[37]) );
  INV_X1 \AddKeyXOR2_XORInst_9_2_U2  ( .A(\AddKeyXOR2_XORInst_9_2_n2 ), .ZN(
        AddRoundKeyOutput[38]) );
  XNOR2_X1 \AddKeyXOR2_XORInst_9_2_U1  ( .A(MCOutput[38]), .B(Key[38]), .ZN(
        \AddKeyXOR2_XORInst_9_2_n2 ) );
  XOR2_X2 \AddKeyXOR2_XORInst_9_3_U1  ( .A(MCOutput[39]), .B(Key[39]), .Z(
        AddRoundKeyOutput[39]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n44 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n43 ), .ZN(
        PermutationInput[0]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n42 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n41 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n40 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n39 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n44 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n38 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n37 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n39 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U20  ( .A1(
        AddRoundKeyOutput[0]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U19  ( .A1(
        CipherErrorVec[2]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n35 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n36 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U18  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n38 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n40 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U16  ( .A1(
        CipherErrorVec[2]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n31 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n32 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U15  ( .A1(
        AddRoundKeyOutput[0]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n31 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n30 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n42 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U12  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n29 ), .B(
        AddRoundKeyOutput[2]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n42 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U11  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n28 ), .A2(
        CipherErrorVec[1]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n29 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U10  ( .A1(
        CipherErrorVec[2]), .A2(CipherErrorVec[0]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U9  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n27 ), .B(
        AddRoundKeyOutput[3]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n26 ), .A2(
        CipherErrorVec[0]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U7  ( .A1(
        CipherErrorVec[2]), .A2(CipherErrorVec[1]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n26 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U6  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n35 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n24 ), .B(
        AddRoundKeyOutput[1]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n33 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U4  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n25 ), .A2(
        CipherErrorVec[2]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U3  ( .A1(
        CipherErrorVec[0]), .A2(CipherErrorVec[1]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n25 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n24 ), .ZN(
        PermutationInput[1]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n23 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n21 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n20 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n22 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U12  ( .A(
        AddRoundKeyOutput[2]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n19 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n23 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U11  ( .A1(
        CipherErrorVec[1]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U10  ( .A1(
        CipherErrorVec[0]), .A2(CipherErrorVec[2]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n18 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U8  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n17 ), .B(
        AddRoundKeyOutput[3]), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n21 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U7  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n16 ), .A2(
        CipherErrorVec[0]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n17 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U6  ( .A(
        AddRoundKeyOutput[0]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n15 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U5  ( .A1(
        CipherErrorVec[0]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n14 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n15 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U4  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n16 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n14 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U3  ( .A1(
        CipherErrorVec[1]), .A2(CipherErrorVec[2]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n16 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U19  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n32 ), .ZN(
        PermutationInput[2]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n29 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n30 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U15  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n25 ), .B(
        AddRoundKeyOutput[2]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n29 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U14  ( .A1(
        CipherErrorVec[1]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n24 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U13  ( .A1(
        CipherErrorVec[2]), .A2(CipherErrorVec[0]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n24 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U12  ( .A(
        AddRoundKeyOutput[1]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n23 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U11  ( .A1(
        CipherErrorVec[2]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n23 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n33 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U9  ( .A(
        AddRoundKeyOutput[0]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n21 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U7  ( .A1(
        CipherErrorVec[1]), .A2(CipherErrorVec[0]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n22 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U6  ( .A(
        CipherErrorVec[2]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n20 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U5  ( .A(
        AddRoundKeyOutput[3]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n19 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n27 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U4  ( .A1(
        CipherErrorVec[0]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U3  ( .A1(
        CipherErrorVec[2]), .A2(CipherErrorVec[1]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n18 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U26  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n48 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n47 ), .ZN(
        PermutationInput[3]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U25  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n46 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n45 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n47 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n44 ), .A2(
        AddRoundKeyOutput[0]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n45 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n43 ), .A2(
        AddRoundKeyOutput[3]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n46 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n42 ), .A2(
        CipherErrorVec[0]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n40 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n48 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U20  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n39 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n38 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n40 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U19  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n44 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n38 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n42 ), .A2(
        AddRoundKeyOutput[3]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n44 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U17  ( .A1(
        CipherErrorVec[0]), .A2(AddRoundKeyOutput[0]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n39 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n37 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n36 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U14  ( .A1(
        CipherErrorVec[0]), .A2(AddRoundKeyOutput[3]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U13  ( .A(
        AddRoundKeyOutput[2]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n33 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n35 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U12  ( .A1(
        CipherErrorVec[1]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n33 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U11  ( .A(
        CipherErrorVec[2]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n29 ), .A2(
        AddRoundKeyOutput[2]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n30 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U8  ( .A1(
        CipherErrorVec[0]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n29 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U7  ( .A(
        AddRoundKeyOutput[3]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n42 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n28 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U6  ( .A1(
        CipherErrorVec[1]), .A2(CipherErrorVec[2]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n42 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n27 ), .B(
        AddRoundKeyOutput[1]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U4  ( .A1(
        CipherErrorVec[2]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U3  ( .A1(
        CipherErrorVec[1]), .A2(CipherErrorVec[0]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n44 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n43 ), .ZN(
        PermutationInput[4]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n42 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n41 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n40 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n39 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n44 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n38 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n37 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n39 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U20  ( .A1(
        AddRoundKeyOutput[4]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U19  ( .A1(
        CipherErrorVec[5]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n35 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n36 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U18  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n38 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n40 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U16  ( .A1(
        CipherErrorVec[5]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n31 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n32 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U15  ( .A1(
        AddRoundKeyOutput[4]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n31 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n30 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n42 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U12  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n29 ), .B(
        AddRoundKeyOutput[6]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n42 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U11  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n28 ), .A2(
        CipherErrorVec[4]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n29 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U10  ( .A1(
        CipherErrorVec[5]), .A2(CipherErrorVec[3]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U9  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n27 ), .B(
        AddRoundKeyOutput[7]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n26 ), .A2(
        CipherErrorVec[3]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U7  ( .A1(
        CipherErrorVec[5]), .A2(CipherErrorVec[4]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n26 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U6  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n35 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n24 ), .B(
        AddRoundKeyOutput[5]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n33 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U4  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n25 ), .A2(
        CipherErrorVec[5]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U3  ( .A1(
        CipherErrorVec[3]), .A2(CipherErrorVec[4]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n25 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n24 ), .ZN(
        PermutationInput[5]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n23 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n21 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n20 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n22 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U12  ( .A(
        AddRoundKeyOutput[6]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n19 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n23 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U11  ( .A1(
        CipherErrorVec[4]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U10  ( .A1(
        CipherErrorVec[3]), .A2(CipherErrorVec[5]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n18 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U8  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n17 ), .B(
        AddRoundKeyOutput[7]), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n21 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U7  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n16 ), .A2(
        CipherErrorVec[3]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n17 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U6  ( .A(
        AddRoundKeyOutput[4]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n15 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U5  ( .A1(
        CipherErrorVec[3]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n14 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n15 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U4  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n16 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n14 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U3  ( .A1(
        CipherErrorVec[4]), .A2(CipherErrorVec[5]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n16 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U19  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n32 ), .ZN(
        PermutationInput[6]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n29 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n30 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U15  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n25 ), .B(
        AddRoundKeyOutput[6]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n29 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U14  ( .A1(
        CipherErrorVec[4]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n24 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U13  ( .A1(
        CipherErrorVec[5]), .A2(CipherErrorVec[3]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n24 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U12  ( .A(
        AddRoundKeyOutput[5]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n23 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U11  ( .A1(
        CipherErrorVec[5]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n23 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n33 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U9  ( .A(
        AddRoundKeyOutput[4]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n21 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U7  ( .A1(
        CipherErrorVec[4]), .A2(CipherErrorVec[3]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n22 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U6  ( .A(
        CipherErrorVec[5]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n20 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U5  ( .A(
        AddRoundKeyOutput[7]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n19 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n27 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U4  ( .A1(
        CipherErrorVec[3]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U3  ( .A1(
        CipherErrorVec[5]), .A2(CipherErrorVec[4]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n18 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U26  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n48 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n47 ), .ZN(
        PermutationInput[7]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U25  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n46 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n45 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n47 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n44 ), .A2(
        AddRoundKeyOutput[4]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n45 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n43 ), .A2(
        AddRoundKeyOutput[7]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n46 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n42 ), .A2(
        CipherErrorVec[3]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n40 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n48 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U20  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n39 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n38 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n40 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U19  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n44 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n38 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n42 ), .A2(
        AddRoundKeyOutput[7]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n44 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U17  ( .A1(
        CipherErrorVec[3]), .A2(AddRoundKeyOutput[4]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n39 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n37 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n36 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U14  ( .A1(
        CipherErrorVec[3]), .A2(AddRoundKeyOutput[7]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U13  ( .A(
        AddRoundKeyOutput[6]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n33 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n35 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U12  ( .A1(
        CipherErrorVec[4]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n33 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U11  ( .A(
        CipherErrorVec[5]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n29 ), .A2(
        AddRoundKeyOutput[6]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n30 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U8  ( .A1(
        CipherErrorVec[3]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n29 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U7  ( .A(
        AddRoundKeyOutput[7]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n42 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n28 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U6  ( .A1(
        CipherErrorVec[4]), .A2(CipherErrorVec[5]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n42 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n27 ), .B(
        AddRoundKeyOutput[5]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U4  ( .A1(
        CipherErrorVec[5]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U3  ( .A1(
        CipherErrorVec[4]), .A2(CipherErrorVec[3]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n44 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n43 ), .ZN(
        PermutationInput[8]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n42 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n41 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n40 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n39 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n44 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n38 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n37 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n39 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U20  ( .A1(
        AddRoundKeyOutput[8]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U19  ( .A1(
        CipherErrorVec[8]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n35 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n36 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U18  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n38 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n40 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U16  ( .A1(
        CipherErrorVec[8]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n31 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n32 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U15  ( .A1(
        AddRoundKeyOutput[8]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n31 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n30 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n42 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U12  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n29 ), .B(
        AddRoundKeyOutput[10]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n42 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U11  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n28 ), .A2(
        CipherErrorVec[7]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n29 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U10  ( .A1(
        CipherErrorVec[8]), .A2(CipherErrorVec[6]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U9  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n27 ), .B(
        AddRoundKeyOutput[11]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n26 ), .A2(
        CipherErrorVec[6]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U7  ( .A1(
        CipherErrorVec[8]), .A2(CipherErrorVec[7]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n26 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U6  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n35 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n24 ), .B(
        AddRoundKeyOutput[9]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n33 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U4  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n25 ), .A2(
        CipherErrorVec[8]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U3  ( .A1(
        CipherErrorVec[6]), .A2(CipherErrorVec[7]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n25 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n24 ), .ZN(
        PermutationInput[9]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n23 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n21 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n20 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n22 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U12  ( .A(
        AddRoundKeyOutput[10]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n19 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n23 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U11  ( .A1(
        CipherErrorVec[7]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U10  ( .A1(
        CipherErrorVec[6]), .A2(CipherErrorVec[8]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n18 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U8  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n17 ), .B(
        AddRoundKeyOutput[11]), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n21 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U7  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n16 ), .A2(
        CipherErrorVec[6]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n17 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U6  ( .A(
        AddRoundKeyOutput[8]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n15 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U5  ( .A1(
        CipherErrorVec[6]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n14 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n15 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U4  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n16 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n14 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U3  ( .A1(
        CipherErrorVec[7]), .A2(CipherErrorVec[8]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n16 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U19  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n32 ), .ZN(
        PermutationInput[10]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n29 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n30 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U15  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n25 ), .B(
        AddRoundKeyOutput[10]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n29 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U14  ( .A1(
        CipherErrorVec[7]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n24 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U13  ( .A1(
        CipherErrorVec[8]), .A2(CipherErrorVec[6]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n24 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U12  ( .A(
        AddRoundKeyOutput[9]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n23 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U11  ( .A1(
        CipherErrorVec[8]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n23 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n33 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U9  ( .A(
        AddRoundKeyOutput[8]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n21 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U7  ( .A1(
        CipherErrorVec[7]), .A2(CipherErrorVec[6]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n22 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U6  ( .A(
        CipherErrorVec[8]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n20 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U5  ( .A(
        AddRoundKeyOutput[11]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n19 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n27 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U4  ( .A1(
        CipherErrorVec[6]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U3  ( .A1(
        CipherErrorVec[8]), .A2(CipherErrorVec[7]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n18 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U26  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n48 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n47 ), .ZN(
        PermutationInput[11]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U25  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n46 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n45 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n47 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n44 ), .A2(
        AddRoundKeyOutput[8]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n45 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n43 ), .A2(
        AddRoundKeyOutput[11]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n46 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n42 ), .A2(
        CipherErrorVec[6]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n40 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n48 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U20  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n39 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n38 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n40 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U19  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n44 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n38 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n42 ), .A2(
        AddRoundKeyOutput[11]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n44 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U17  ( .A1(
        CipherErrorVec[6]), .A2(AddRoundKeyOutput[8]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n39 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n37 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n36 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U14  ( .A1(
        CipherErrorVec[6]), .A2(AddRoundKeyOutput[11]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U13  ( .A(
        AddRoundKeyOutput[10]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n33 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n35 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U12  ( .A1(
        CipherErrorVec[7]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n33 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U11  ( .A(
        CipherErrorVec[8]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n29 ), .A2(
        AddRoundKeyOutput[10]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n30 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U8  ( .A1(
        CipherErrorVec[6]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n29 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U7  ( .A(
        AddRoundKeyOutput[11]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n42 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n28 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U6  ( .A1(
        CipherErrorVec[7]), .A2(CipherErrorVec[8]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n42 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n27 ), .B(
        AddRoundKeyOutput[9]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U4  ( .A1(
        CipherErrorVec[8]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U3  ( .A1(
        CipherErrorVec[7]), .A2(CipherErrorVec[6]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n44 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n43 ), .ZN(
        PermutationInput[12]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n42 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n41 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n40 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n39 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n44 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n38 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n37 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n39 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U20  ( .A1(
        AddRoundKeyOutput[12]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U19  ( .A1(
        CipherErrorVec[11]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n35 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n36 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U18  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n38 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n40 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U16  ( .A1(
        CipherErrorVec[11]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n31 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n32 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U15  ( .A1(
        AddRoundKeyOutput[12]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n31 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n30 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n42 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U12  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n29 ), .B(
        AddRoundKeyOutput[14]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n42 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U11  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n28 ), .A2(
        CipherErrorVec[10]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n29 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U10  ( .A1(
        CipherErrorVec[11]), .A2(CipherErrorVec[9]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U9  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n27 ), .B(
        AddRoundKeyOutput[15]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n26 ), .A2(
        CipherErrorVec[9]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U7  ( .A1(
        CipherErrorVec[11]), .A2(CipherErrorVec[10]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n26 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U6  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n35 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n24 ), .B(
        AddRoundKeyOutput[13]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n33 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U4  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n25 ), .A2(
        CipherErrorVec[11]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U3  ( .A1(
        CipherErrorVec[9]), .A2(CipherErrorVec[10]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n25 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n24 ), .ZN(
        PermutationInput[13]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n23 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n21 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n20 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n22 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U12  ( .A(
        AddRoundKeyOutput[14]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n19 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n23 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U11  ( .A1(
        CipherErrorVec[10]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U10  ( .A1(
        CipherErrorVec[9]), .A2(CipherErrorVec[11]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n18 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U8  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n17 ), .B(
        AddRoundKeyOutput[15]), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n21 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U7  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n16 ), .A2(
        CipherErrorVec[9]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n17 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U6  ( .A(
        AddRoundKeyOutput[12]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n15 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U5  ( .A1(
        CipherErrorVec[9]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n14 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n15 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U4  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n16 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n14 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U3  ( .A1(
        CipherErrorVec[10]), .A2(CipherErrorVec[11]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n16 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U19  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n32 ), .ZN(
        PermutationInput[14]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n29 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n30 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U15  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n25 ), .B(
        AddRoundKeyOutput[14]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n29 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U14  ( .A1(
        CipherErrorVec[10]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n24 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U13  ( .A1(
        CipherErrorVec[11]), .A2(CipherErrorVec[9]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n24 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U12  ( .A(
        AddRoundKeyOutput[13]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n23 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U11  ( .A1(
        CipherErrorVec[11]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n23 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n33 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U9  ( .A(
        AddRoundKeyOutput[12]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n21 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U7  ( .A1(
        CipherErrorVec[10]), .A2(CipherErrorVec[9]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n22 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U6  ( .A(
        CipherErrorVec[11]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n20 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U5  ( .A(
        AddRoundKeyOutput[15]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n19 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n27 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U4  ( .A1(
        CipherErrorVec[9]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U3  ( .A1(
        CipherErrorVec[11]), .A2(CipherErrorVec[10]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n18 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U26  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n48 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n47 ), .ZN(
        PermutationInput[15]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U25  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n46 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n45 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n47 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n44 ), .A2(
        AddRoundKeyOutput[12]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n45 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n43 ), .A2(
        AddRoundKeyOutput[15]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n46 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n42 ), .A2(
        CipherErrorVec[9]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n40 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n48 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U20  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n39 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n38 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n40 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U19  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n44 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n38 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n42 ), .A2(
        AddRoundKeyOutput[15]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n44 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U17  ( .A1(
        CipherErrorVec[9]), .A2(AddRoundKeyOutput[12]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n39 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n37 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n36 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U14  ( .A1(
        CipherErrorVec[9]), .A2(AddRoundKeyOutput[15]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U13  ( .A(
        AddRoundKeyOutput[14]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n33 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n35 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U12  ( .A1(
        CipherErrorVec[10]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n33 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U11  ( .A(
        CipherErrorVec[11]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n29 ), .A2(
        AddRoundKeyOutput[14]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n30 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U8  ( .A1(
        CipherErrorVec[9]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n29 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U7  ( .A(
        AddRoundKeyOutput[15]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n42 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n28 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U6  ( .A1(
        CipherErrorVec[10]), .A2(CipherErrorVec[11]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n42 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n27 ), .B(
        AddRoundKeyOutput[13]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U4  ( .A1(
        CipherErrorVec[11]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U3  ( .A1(
        CipherErrorVec[10]), .A2(CipherErrorVec[9]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n44 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n43 ), .ZN(
        PermutationInput[16]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n42 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n41 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n40 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n39 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n44 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n38 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n37 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n39 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U20  ( .A1(
        AddRoundKeyOutput[16]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U19  ( .A1(
        CipherErrorVec[14]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n35 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n36 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U18  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n38 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n40 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U16  ( .A1(
        CipherErrorVec[14]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n31 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n32 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U15  ( .A1(
        AddRoundKeyOutput[16]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n31 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n30 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n42 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U12  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n29 ), .B(
        AddRoundKeyOutput[18]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n42 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U11  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n28 ), .A2(
        CipherErrorVec[13]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n29 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U10  ( .A1(
        CipherErrorVec[14]), .A2(CipherErrorVec[12]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U9  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n27 ), .B(
        AddRoundKeyOutput[19]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n26 ), .A2(
        CipherErrorVec[12]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U7  ( .A1(
        CipherErrorVec[14]), .A2(CipherErrorVec[13]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n26 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U6  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n35 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n24 ), .B(
        AddRoundKeyOutput[17]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n33 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U4  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n25 ), .A2(
        CipherErrorVec[14]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U3  ( .A1(
        CipherErrorVec[12]), .A2(CipherErrorVec[13]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n25 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n24 ), .ZN(
        PermutationInput[17]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n23 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n21 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n20 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n22 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U12  ( .A(
        AddRoundKeyOutput[18]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n19 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n23 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U11  ( .A1(
        CipherErrorVec[13]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U10  ( .A1(
        CipherErrorVec[12]), .A2(CipherErrorVec[14]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n18 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U8  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n17 ), .B(
        AddRoundKeyOutput[19]), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n21 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U7  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n16 ), .A2(
        CipherErrorVec[12]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n17 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U6  ( .A(
        AddRoundKeyOutput[16]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n15 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U5  ( .A1(
        CipherErrorVec[12]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n14 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n15 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U4  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n16 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n14 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U3  ( .A1(
        CipherErrorVec[13]), .A2(CipherErrorVec[14]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n16 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U19  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n32 ), .ZN(
        PermutationInput[18]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n29 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n30 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U15  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n25 ), .B(
        AddRoundKeyOutput[18]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n29 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U14  ( .A1(
        CipherErrorVec[13]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n24 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U13  ( .A1(
        CipherErrorVec[14]), .A2(CipherErrorVec[12]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n24 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U12  ( .A(
        AddRoundKeyOutput[17]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n23 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U11  ( .A1(
        CipherErrorVec[14]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n23 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n33 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U9  ( .A(
        AddRoundKeyOutput[16]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n21 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U7  ( .A1(
        CipherErrorVec[13]), .A2(CipherErrorVec[12]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n22 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U6  ( .A(
        CipherErrorVec[14]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n20 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U5  ( .A(
        AddRoundKeyOutput[19]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n19 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n27 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U4  ( .A1(
        CipherErrorVec[12]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U3  ( .A1(
        CipherErrorVec[14]), .A2(CipherErrorVec[13]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n18 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U26  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n48 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n47 ), .ZN(
        PermutationInput[19]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U25  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n46 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n45 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n47 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n44 ), .A2(
        AddRoundKeyOutput[16]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n45 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n43 ), .A2(
        AddRoundKeyOutput[19]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n46 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n42 ), .A2(
        CipherErrorVec[12]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n40 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n48 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U20  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n39 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n38 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n40 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U19  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n44 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n38 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n42 ), .A2(
        AddRoundKeyOutput[19]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n44 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U17  ( .A1(
        CipherErrorVec[12]), .A2(AddRoundKeyOutput[16]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n39 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n37 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n36 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U14  ( .A1(
        CipherErrorVec[12]), .A2(AddRoundKeyOutput[19]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U13  ( .A(
        AddRoundKeyOutput[18]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n33 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n35 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U12  ( .A1(
        CipherErrorVec[13]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n33 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U11  ( .A(
        CipherErrorVec[14]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n29 ), .A2(
        AddRoundKeyOutput[18]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n30 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U8  ( .A1(
        CipherErrorVec[12]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n29 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U7  ( .A(
        AddRoundKeyOutput[19]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n42 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n28 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U6  ( .A1(
        CipherErrorVec[13]), .A2(CipherErrorVec[14]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n42 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n27 ), .B(
        AddRoundKeyOutput[17]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U4  ( .A1(
        CipherErrorVec[14]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U3  ( .A1(
        CipherErrorVec[13]), .A2(CipherErrorVec[12]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n44 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n43 ), .ZN(
        PermutationInput[20]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n42 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n41 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n40 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n39 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n44 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n38 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n37 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n39 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U20  ( .A1(
        AddRoundKeyOutput[20]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U19  ( .A1(
        CipherErrorVec[17]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n35 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n36 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U18  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n38 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n40 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U16  ( .A1(
        CipherErrorVec[17]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n31 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n32 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U15  ( .A1(
        AddRoundKeyOutput[20]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n31 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n30 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n42 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U12  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n29 ), .B(
        AddRoundKeyOutput[22]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n42 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U11  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n28 ), .A2(
        CipherErrorVec[16]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n29 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U10  ( .A1(
        CipherErrorVec[17]), .A2(CipherErrorVec[15]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U9  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n27 ), .B(
        AddRoundKeyOutput[23]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n26 ), .A2(
        CipherErrorVec[15]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U7  ( .A1(
        CipherErrorVec[17]), .A2(CipherErrorVec[16]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n26 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U6  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n35 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n24 ), .B(
        AddRoundKeyOutput[21]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n33 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U4  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n25 ), .A2(
        CipherErrorVec[17]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U3  ( .A1(
        CipherErrorVec[15]), .A2(CipherErrorVec[16]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n25 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n24 ), .ZN(
        PermutationInput[21]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n23 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n21 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n20 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n22 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U12  ( .A(
        AddRoundKeyOutput[22]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n19 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n23 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U11  ( .A1(
        CipherErrorVec[16]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U10  ( .A1(
        CipherErrorVec[15]), .A2(CipherErrorVec[17]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n18 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U8  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n17 ), .B(
        AddRoundKeyOutput[23]), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n21 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U7  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n16 ), .A2(
        CipherErrorVec[15]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n17 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U6  ( .A(
        AddRoundKeyOutput[20]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n15 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U5  ( .A1(
        CipherErrorVec[15]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n14 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n15 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U4  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n16 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n14 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U3  ( .A1(
        CipherErrorVec[16]), .A2(CipherErrorVec[17]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n16 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U19  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n32 ), .ZN(
        PermutationInput[22]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n29 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n30 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U15  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n25 ), .B(
        AddRoundKeyOutput[22]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n29 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U14  ( .A1(
        CipherErrorVec[16]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n24 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U13  ( .A1(
        CipherErrorVec[17]), .A2(CipherErrorVec[15]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n24 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U12  ( .A(
        AddRoundKeyOutput[21]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n23 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U11  ( .A1(
        CipherErrorVec[17]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n23 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n33 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U9  ( .A(
        AddRoundKeyOutput[20]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n21 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U7  ( .A1(
        CipherErrorVec[16]), .A2(CipherErrorVec[15]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n22 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U6  ( .A(
        CipherErrorVec[17]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n20 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U5  ( .A(
        AddRoundKeyOutput[23]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n19 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n27 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U4  ( .A1(
        CipherErrorVec[15]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U3  ( .A1(
        CipherErrorVec[17]), .A2(CipherErrorVec[16]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n18 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U26  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n48 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n47 ), .ZN(
        PermutationInput[23]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U25  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n46 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n45 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n47 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n44 ), .A2(
        AddRoundKeyOutput[20]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n45 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n43 ), .A2(
        AddRoundKeyOutput[23]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n46 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n42 ), .A2(
        CipherErrorVec[15]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n40 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n48 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U20  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n39 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n38 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n40 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U19  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n44 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n38 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n42 ), .A2(
        AddRoundKeyOutput[23]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n44 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U17  ( .A1(
        CipherErrorVec[15]), .A2(AddRoundKeyOutput[20]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n39 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n37 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n36 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U14  ( .A1(
        CipherErrorVec[15]), .A2(AddRoundKeyOutput[23]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U13  ( .A(
        AddRoundKeyOutput[22]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n33 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n35 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U12  ( .A1(
        CipherErrorVec[16]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n33 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U11  ( .A(
        CipherErrorVec[17]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n29 ), .A2(
        AddRoundKeyOutput[22]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n30 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U8  ( .A1(
        CipherErrorVec[15]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n29 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U7  ( .A(
        AddRoundKeyOutput[23]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n42 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n28 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U6  ( .A1(
        CipherErrorVec[16]), .A2(CipherErrorVec[17]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n42 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n27 ), .B(
        AddRoundKeyOutput[21]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U4  ( .A1(
        CipherErrorVec[17]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U3  ( .A1(
        CipherErrorVec[16]), .A2(CipherErrorVec[15]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n44 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n43 ), .ZN(
        PermutationInput[24]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n42 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n41 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n40 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n39 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n44 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n38 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n37 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n39 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U20  ( .A1(
        AddRoundKeyOutput[24]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U19  ( .A1(
        CipherErrorVec[20]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n35 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n36 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U18  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n38 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n40 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U16  ( .A1(
        CipherErrorVec[20]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n31 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n32 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U15  ( .A1(
        AddRoundKeyOutput[24]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n31 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n30 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n42 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U12  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n29 ), .B(
        AddRoundKeyOutput[26]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n42 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U11  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n28 ), .A2(
        CipherErrorVec[19]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n29 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U10  ( .A1(
        CipherErrorVec[20]), .A2(CipherErrorVec[18]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U9  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n27 ), .B(
        AddRoundKeyOutput[27]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n26 ), .A2(
        CipherErrorVec[18]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U7  ( .A1(
        CipherErrorVec[20]), .A2(CipherErrorVec[19]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n26 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U6  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n35 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n24 ), .B(
        AddRoundKeyOutput[25]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n33 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U4  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n25 ), .A2(
        CipherErrorVec[20]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U3  ( .A1(
        CipherErrorVec[18]), .A2(CipherErrorVec[19]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n25 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n24 ), .ZN(
        PermutationInput[25]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n23 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n21 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n20 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n22 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U12  ( .A(
        AddRoundKeyOutput[26]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n19 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n23 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U11  ( .A1(
        CipherErrorVec[19]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U10  ( .A1(
        CipherErrorVec[18]), .A2(CipherErrorVec[20]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n18 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U8  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n17 ), .B(
        AddRoundKeyOutput[27]), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n21 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U7  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n16 ), .A2(
        CipherErrorVec[18]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n17 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U6  ( .A(
        AddRoundKeyOutput[24]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n15 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U5  ( .A1(
        CipherErrorVec[18]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n14 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n15 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U4  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n16 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n14 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U3  ( .A1(
        CipherErrorVec[19]), .A2(CipherErrorVec[20]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n16 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U19  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n32 ), .ZN(
        PermutationInput[26]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n29 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n30 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U15  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n25 ), .B(
        AddRoundKeyOutput[26]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n29 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U14  ( .A1(
        CipherErrorVec[19]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n24 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U13  ( .A1(
        CipherErrorVec[20]), .A2(CipherErrorVec[18]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n24 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U12  ( .A(
        AddRoundKeyOutput[25]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n23 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U11  ( .A1(
        CipherErrorVec[20]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n23 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n33 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U9  ( .A(
        AddRoundKeyOutput[24]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n21 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U7  ( .A1(
        CipherErrorVec[19]), .A2(CipherErrorVec[18]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n22 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U6  ( .A(
        CipherErrorVec[20]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n20 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U5  ( .A(
        AddRoundKeyOutput[27]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n19 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n27 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U4  ( .A1(
        CipherErrorVec[18]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U3  ( .A1(
        CipherErrorVec[20]), .A2(CipherErrorVec[19]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n18 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U26  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n48 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n47 ), .ZN(
        PermutationInput[27]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U25  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n46 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n45 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n47 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n44 ), .A2(
        AddRoundKeyOutput[24]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n45 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n43 ), .A2(
        AddRoundKeyOutput[27]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n46 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n42 ), .A2(
        CipherErrorVec[18]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n40 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n48 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U20  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n39 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n38 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n40 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U19  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n44 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n38 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n42 ), .A2(
        AddRoundKeyOutput[27]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n44 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U17  ( .A1(
        CipherErrorVec[18]), .A2(AddRoundKeyOutput[24]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n39 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n37 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n36 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U14  ( .A1(
        CipherErrorVec[18]), .A2(AddRoundKeyOutput[27]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U13  ( .A(
        AddRoundKeyOutput[26]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n33 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n35 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U12  ( .A1(
        CipherErrorVec[19]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n33 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U11  ( .A(
        CipherErrorVec[20]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n29 ), .A2(
        AddRoundKeyOutput[26]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n30 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U8  ( .A1(
        CipherErrorVec[18]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n29 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U7  ( .A(
        AddRoundKeyOutput[27]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n42 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n28 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U6  ( .A1(
        CipherErrorVec[19]), .A2(CipherErrorVec[20]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n42 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n27 ), .B(
        AddRoundKeyOutput[25]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U4  ( .A1(
        CipherErrorVec[20]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U3  ( .A1(
        CipherErrorVec[19]), .A2(CipherErrorVec[18]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n44 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n43 ), .ZN(
        PermutationInput[28]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n42 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n41 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n40 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n39 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n44 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n38 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n37 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n39 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U20  ( .A1(
        AddRoundKeyOutput[28]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U19  ( .A1(
        CipherErrorVec[23]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n35 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n36 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U18  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n38 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n40 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U16  ( .A1(
        CipherErrorVec[23]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n31 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n32 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U15  ( .A1(
        AddRoundKeyOutput[28]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n31 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n30 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n42 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U12  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n29 ), .B(
        AddRoundKeyOutput[30]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n42 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U11  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n28 ), .A2(
        CipherErrorVec[22]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n29 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U10  ( .A1(
        CipherErrorVec[23]), .A2(CipherErrorVec[21]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U9  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n27 ), .B(
        AddRoundKeyOutput[31]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n26 ), .A2(
        CipherErrorVec[21]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U7  ( .A1(
        CipherErrorVec[23]), .A2(CipherErrorVec[22]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n26 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U6  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n35 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n24 ), .B(
        AddRoundKeyOutput[29]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n33 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U4  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n25 ), .A2(
        CipherErrorVec[23]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U3  ( .A1(
        CipherErrorVec[21]), .A2(CipherErrorVec[22]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n25 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n24 ), .ZN(
        PermutationInput[29]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n23 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n21 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n20 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n22 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U12  ( .A(
        AddRoundKeyOutput[30]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n19 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n23 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U11  ( .A1(
        CipherErrorVec[22]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U10  ( .A1(
        CipherErrorVec[21]), .A2(CipherErrorVec[23]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n18 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U8  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n17 ), .B(
        AddRoundKeyOutput[31]), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n21 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U7  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n16 ), .A2(
        CipherErrorVec[21]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n17 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U6  ( .A(
        AddRoundKeyOutput[28]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n15 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U5  ( .A1(
        CipherErrorVec[21]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n14 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n15 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U4  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n16 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n14 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U3  ( .A1(
        CipherErrorVec[22]), .A2(CipherErrorVec[23]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n16 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U19  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n32 ), .ZN(
        PermutationInput[30]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n29 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n30 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U15  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n25 ), .B(
        AddRoundKeyOutput[30]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n29 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U14  ( .A1(
        CipherErrorVec[22]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n24 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U13  ( .A1(
        CipherErrorVec[23]), .A2(CipherErrorVec[21]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n24 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U12  ( .A(
        AddRoundKeyOutput[29]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n23 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U11  ( .A1(
        CipherErrorVec[23]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n23 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n33 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U9  ( .A(
        AddRoundKeyOutput[28]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n21 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U7  ( .A1(
        CipherErrorVec[22]), .A2(CipherErrorVec[21]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n22 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U6  ( .A(
        CipherErrorVec[23]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n20 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U5  ( .A(
        AddRoundKeyOutput[31]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n19 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n27 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U4  ( .A1(
        CipherErrorVec[21]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U3  ( .A1(
        CipherErrorVec[23]), .A2(CipherErrorVec[22]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n18 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U26  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n48 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n47 ), .ZN(
        PermutationInput[31]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U25  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n46 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n45 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n47 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n44 ), .A2(
        AddRoundKeyOutput[28]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n45 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n43 ), .A2(
        AddRoundKeyOutput[31]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n46 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n42 ), .A2(
        CipherErrorVec[21]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n40 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n48 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U20  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n39 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n38 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n40 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U19  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n44 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n38 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n42 ), .A2(
        AddRoundKeyOutput[31]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n44 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U17  ( .A1(
        CipherErrorVec[21]), .A2(AddRoundKeyOutput[28]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n39 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n37 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n36 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U14  ( .A1(
        CipherErrorVec[21]), .A2(AddRoundKeyOutput[31]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U13  ( .A(
        AddRoundKeyOutput[30]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n33 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n35 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U12  ( .A1(
        CipherErrorVec[22]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n33 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U11  ( .A(
        CipherErrorVec[23]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n29 ), .A2(
        AddRoundKeyOutput[30]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n30 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U8  ( .A1(
        CipherErrorVec[21]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n29 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U7  ( .A(
        AddRoundKeyOutput[31]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n42 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n28 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U6  ( .A1(
        CipherErrorVec[22]), .A2(CipherErrorVec[23]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n42 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n27 ), .B(
        AddRoundKeyOutput[29]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U4  ( .A1(
        CipherErrorVec[23]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U3  ( .A1(
        CipherErrorVec[22]), .A2(CipherErrorVec[21]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n44 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n43 ), .ZN(
        PermutationInput[32]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n42 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n41 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n40 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n39 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n44 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n38 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n37 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n39 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U20  ( .A1(
        AddRoundKeyOutput[32]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U19  ( .A1(
        CipherErrorVec[26]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n35 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n36 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U18  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n38 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n40 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U16  ( .A1(
        CipherErrorVec[26]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n31 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n32 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U15  ( .A1(
        AddRoundKeyOutput[32]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n31 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n30 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n42 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U12  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n29 ), .B(
        AddRoundKeyOutput[34]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n42 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U11  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n28 ), .A2(
        CipherErrorVec[25]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n29 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U10  ( .A1(
        CipherErrorVec[26]), .A2(CipherErrorVec[24]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U9  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n27 ), .B(
        AddRoundKeyOutput[35]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n26 ), .A2(
        CipherErrorVec[24]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U7  ( .A1(
        CipherErrorVec[26]), .A2(CipherErrorVec[25]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n26 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U6  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n35 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n24 ), .B(
        AddRoundKeyOutput[33]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n33 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U4  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n25 ), .A2(
        CipherErrorVec[26]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U3  ( .A1(
        CipherErrorVec[24]), .A2(CipherErrorVec[25]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n25 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n24 ), .ZN(
        PermutationInput[33]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n23 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n21 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n20 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n22 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U12  ( .A(
        AddRoundKeyOutput[34]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n19 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n23 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U11  ( .A1(
        CipherErrorVec[25]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U10  ( .A1(
        CipherErrorVec[24]), .A2(CipherErrorVec[26]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n18 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U8  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n17 ), .B(
        AddRoundKeyOutput[35]), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n21 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U7  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n16 ), .A2(
        CipherErrorVec[24]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n17 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U6  ( .A(
        AddRoundKeyOutput[32]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n15 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U5  ( .A1(
        CipherErrorVec[24]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n14 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n15 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U4  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n16 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n14 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U3  ( .A1(
        CipherErrorVec[25]), .A2(CipherErrorVec[26]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n16 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U19  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n32 ), .ZN(
        PermutationInput[34]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n29 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n30 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U15  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n25 ), .B(
        AddRoundKeyOutput[34]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n29 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U14  ( .A1(
        CipherErrorVec[25]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n24 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U13  ( .A1(
        CipherErrorVec[26]), .A2(CipherErrorVec[24]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n24 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U12  ( .A(
        AddRoundKeyOutput[33]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n23 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U11  ( .A1(
        CipherErrorVec[26]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n23 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n33 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U9  ( .A(
        AddRoundKeyOutput[32]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n21 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U7  ( .A1(
        CipherErrorVec[25]), .A2(CipherErrorVec[24]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n22 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U6  ( .A(
        CipherErrorVec[26]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n20 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U5  ( .A(
        AddRoundKeyOutput[35]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n19 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n27 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U4  ( .A1(
        CipherErrorVec[24]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U3  ( .A1(
        CipherErrorVec[26]), .A2(CipherErrorVec[25]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n18 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U26  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n48 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n47 ), .ZN(
        PermutationInput[35]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U25  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n46 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n45 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n47 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n44 ), .A2(
        AddRoundKeyOutput[32]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n45 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n43 ), .A2(
        AddRoundKeyOutput[35]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n46 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n42 ), .A2(
        CipherErrorVec[24]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n40 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n48 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U20  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n39 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n38 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n40 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U19  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n44 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n38 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n42 ), .A2(
        AddRoundKeyOutput[35]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n44 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U17  ( .A1(
        CipherErrorVec[24]), .A2(AddRoundKeyOutput[32]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n39 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n37 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n36 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U14  ( .A1(
        CipherErrorVec[24]), .A2(AddRoundKeyOutput[35]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U13  ( .A(
        AddRoundKeyOutput[34]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n33 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n35 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U12  ( .A1(
        CipherErrorVec[25]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n33 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U11  ( .A(
        CipherErrorVec[26]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n29 ), .A2(
        AddRoundKeyOutput[34]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n30 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U8  ( .A1(
        CipherErrorVec[24]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n29 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U7  ( .A(
        AddRoundKeyOutput[35]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n42 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n28 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U6  ( .A1(
        CipherErrorVec[25]), .A2(CipherErrorVec[26]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n42 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n27 ), .B(
        AddRoundKeyOutput[33]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U4  ( .A1(
        CipherErrorVec[26]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U3  ( .A1(
        CipherErrorVec[25]), .A2(CipherErrorVec[24]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n44 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n43 ), .ZN(
        PermutationInput[36]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n42 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n41 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n40 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n39 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n44 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n38 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n37 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n39 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U20  ( .A1(
        AddRoundKeyOutput[36]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U19  ( .A1(
        CipherErrorVec[29]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n35 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n36 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U18  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n38 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n40 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U16  ( .A1(
        CipherErrorVec[29]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n31 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n32 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U15  ( .A1(
        AddRoundKeyOutput[36]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n31 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n30 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n42 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U12  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n29 ), .B(
        AddRoundKeyOutput[38]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n42 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U11  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n28 ), .A2(
        CipherErrorVec[28]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n29 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U10  ( .A1(
        CipherErrorVec[29]), .A2(CipherErrorVec[27]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U9  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n27 ), .B(
        AddRoundKeyOutput[39]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n26 ), .A2(
        CipherErrorVec[27]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U7  ( .A1(
        CipherErrorVec[29]), .A2(CipherErrorVec[28]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n26 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U6  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n35 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n24 ), .B(
        AddRoundKeyOutput[37]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n33 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U4  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n25 ), .A2(
        CipherErrorVec[29]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U3  ( .A1(
        CipherErrorVec[27]), .A2(CipherErrorVec[28]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n25 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n24 ), .ZN(
        PermutationInput[37]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n23 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n21 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n20 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n22 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U12  ( .A(
        AddRoundKeyOutput[38]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n19 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n23 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U11  ( .A1(
        CipherErrorVec[28]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U10  ( .A1(
        CipherErrorVec[27]), .A2(CipherErrorVec[29]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n18 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U8  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n17 ), .B(
        AddRoundKeyOutput[39]), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n21 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U7  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n16 ), .A2(
        CipherErrorVec[27]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n17 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U6  ( .A(
        AddRoundKeyOutput[36]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n15 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U5  ( .A1(
        CipherErrorVec[27]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n14 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n15 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U4  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n16 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n14 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U3  ( .A1(
        CipherErrorVec[28]), .A2(CipherErrorVec[29]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n16 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U19  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n32 ), .ZN(
        PermutationInput[38]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n29 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n30 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U15  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n25 ), .B(
        AddRoundKeyOutput[38]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n29 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U14  ( .A1(
        CipherErrorVec[28]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n24 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U13  ( .A1(
        CipherErrorVec[29]), .A2(CipherErrorVec[27]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n24 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U12  ( .A(
        AddRoundKeyOutput[37]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n23 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U11  ( .A1(
        CipherErrorVec[29]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n23 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n33 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U9  ( .A(
        AddRoundKeyOutput[36]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n21 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U7  ( .A1(
        CipherErrorVec[28]), .A2(CipherErrorVec[27]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n22 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U6  ( .A(
        CipherErrorVec[29]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n20 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U5  ( .A(
        AddRoundKeyOutput[39]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n19 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n27 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U4  ( .A1(
        CipherErrorVec[27]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U3  ( .A1(
        CipherErrorVec[29]), .A2(CipherErrorVec[28]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n18 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U26  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n48 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n47 ), .ZN(
        PermutationInput[39]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U25  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n46 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n45 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n47 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n44 ), .A2(
        AddRoundKeyOutput[36]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n45 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n43 ), .A2(
        AddRoundKeyOutput[39]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n46 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n42 ), .A2(
        CipherErrorVec[27]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n40 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n48 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U20  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n39 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n38 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n40 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U19  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n44 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n38 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n42 ), .A2(
        AddRoundKeyOutput[39]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n44 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U17  ( .A1(
        CipherErrorVec[27]), .A2(AddRoundKeyOutput[36]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n39 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n37 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n36 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U14  ( .A1(
        CipherErrorVec[27]), .A2(AddRoundKeyOutput[39]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U13  ( .A(
        AddRoundKeyOutput[38]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n33 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n35 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U12  ( .A1(
        CipherErrorVec[28]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n33 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U11  ( .A(
        CipherErrorVec[29]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n29 ), .A2(
        AddRoundKeyOutput[38]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n30 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U8  ( .A1(
        CipherErrorVec[27]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n29 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U7  ( .A(
        AddRoundKeyOutput[39]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n42 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n28 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U6  ( .A1(
        CipherErrorVec[28]), .A2(CipherErrorVec[29]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n42 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n27 ), .B(
        AddRoundKeyOutput[37]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U4  ( .A1(
        CipherErrorVec[29]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U3  ( .A1(
        CipherErrorVec[28]), .A2(CipherErrorVec[27]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n44 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n43 ), .ZN(
        PermutationInput[40]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n42 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n41 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n40 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n39 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n44 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n38 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n37 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n39 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U20  ( .A1(
        AddRoundKeyOutput[40]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U19  ( .A1(
        CipherErrorVec[32]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n35 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n36 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U18  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n38 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n40 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U16  ( .A1(
        CipherErrorVec[32]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n31 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n32 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U15  ( .A1(
        AddRoundKeyOutput[40]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n31 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n30 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n42 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U12  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n29 ), .B(
        AddRoundKeyOutput[42]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n42 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U11  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n28 ), .A2(
        CipherErrorVec[31]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n29 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U10  ( .A1(
        CipherErrorVec[32]), .A2(CipherErrorVec[30]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U9  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n27 ), .B(
        AddRoundKeyOutput[43]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n26 ), .A2(
        CipherErrorVec[30]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U7  ( .A1(
        CipherErrorVec[32]), .A2(CipherErrorVec[31]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n26 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U6  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n35 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n24 ), .B(
        AddRoundKeyOutput[41]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n33 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U4  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n25 ), .A2(
        CipherErrorVec[32]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U3  ( .A1(
        CipherErrorVec[30]), .A2(CipherErrorVec[31]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n25 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n24 ), .ZN(
        PermutationInput[41]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n23 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n21 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n20 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n22 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U12  ( .A(
        AddRoundKeyOutput[42]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n19 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n23 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U11  ( .A1(
        CipherErrorVec[31]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U10  ( .A1(
        CipherErrorVec[30]), .A2(CipherErrorVec[32]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n18 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U8  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n17 ), .B(
        AddRoundKeyOutput[43]), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n21 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U7  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n16 ), .A2(
        CipherErrorVec[30]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n17 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U6  ( .A(
        AddRoundKeyOutput[40]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n15 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U5  ( .A1(
        CipherErrorVec[30]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n14 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n15 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U4  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n16 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n14 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U3  ( .A1(
        CipherErrorVec[31]), .A2(CipherErrorVec[32]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n16 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U19  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n32 ), .ZN(
        PermutationInput[42]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n29 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n30 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U15  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n25 ), .B(
        AddRoundKeyOutput[42]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n29 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U14  ( .A1(
        CipherErrorVec[31]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n24 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U13  ( .A1(
        CipherErrorVec[32]), .A2(CipherErrorVec[30]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n24 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U12  ( .A(
        AddRoundKeyOutput[41]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n23 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U11  ( .A1(
        CipherErrorVec[32]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n23 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n33 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U9  ( .A(
        AddRoundKeyOutput[40]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n21 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U7  ( .A1(
        CipherErrorVec[31]), .A2(CipherErrorVec[30]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n22 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U6  ( .A(
        CipherErrorVec[32]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n20 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U5  ( .A(
        AddRoundKeyOutput[43]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n19 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n27 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U4  ( .A1(
        CipherErrorVec[30]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U3  ( .A1(
        CipherErrorVec[32]), .A2(CipherErrorVec[31]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n18 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U26  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n48 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n47 ), .ZN(
        PermutationInput[43]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U25  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n46 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n45 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n47 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n44 ), .A2(
        AddRoundKeyOutput[40]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n45 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n43 ), .A2(
        AddRoundKeyOutput[43]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n46 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n42 ), .A2(
        CipherErrorVec[30]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n40 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n48 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U20  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n39 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n38 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n40 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U19  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n44 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n38 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n42 ), .A2(
        AddRoundKeyOutput[43]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n44 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U17  ( .A1(
        CipherErrorVec[30]), .A2(AddRoundKeyOutput[40]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n39 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n37 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n36 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U14  ( .A1(
        CipherErrorVec[30]), .A2(AddRoundKeyOutput[43]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U13  ( .A(
        AddRoundKeyOutput[42]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n33 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n35 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U12  ( .A1(
        CipherErrorVec[31]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n33 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U11  ( .A(
        CipherErrorVec[32]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n29 ), .A2(
        AddRoundKeyOutput[42]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n30 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U8  ( .A1(
        CipherErrorVec[30]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n29 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U7  ( .A(
        AddRoundKeyOutput[43]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n42 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n28 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U6  ( .A1(
        CipherErrorVec[31]), .A2(CipherErrorVec[32]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n42 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n27 ), .B(
        AddRoundKeyOutput[41]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U4  ( .A1(
        CipherErrorVec[32]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U3  ( .A1(
        CipherErrorVec[31]), .A2(CipherErrorVec[30]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n44 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n43 ), .ZN(
        PermutationInput[44]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n42 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n41 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n40 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n39 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n44 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n38 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n37 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n39 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U20  ( .A1(
        AddRoundKeyOutput[44]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U19  ( .A1(
        CipherErrorVec[35]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n35 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n36 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U18  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n38 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n40 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U16  ( .A1(
        CipherErrorVec[35]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n31 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n32 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U15  ( .A1(
        AddRoundKeyOutput[44]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n31 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n30 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n42 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U12  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n29 ), .B(
        AddRoundKeyOutput[46]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n42 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U11  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n28 ), .A2(
        CipherErrorVec[34]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n29 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U10  ( .A1(
        CipherErrorVec[35]), .A2(CipherErrorVec[33]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U9  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n27 ), .B(
        AddRoundKeyOutput[47]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n26 ), .A2(
        CipherErrorVec[33]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U7  ( .A1(
        CipherErrorVec[35]), .A2(CipherErrorVec[34]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n26 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U6  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n35 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n24 ), .B(
        AddRoundKeyOutput[45]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n33 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U4  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n25 ), .A2(
        CipherErrorVec[35]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U3  ( .A1(
        CipherErrorVec[33]), .A2(CipherErrorVec[34]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n25 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n24 ), .ZN(
        PermutationInput[45]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n23 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n21 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n20 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n22 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U12  ( .A(
        AddRoundKeyOutput[46]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n19 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n23 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U11  ( .A1(
        CipherErrorVec[34]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U10  ( .A1(
        CipherErrorVec[33]), .A2(CipherErrorVec[35]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n18 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U8  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n17 ), .B(
        AddRoundKeyOutput[47]), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n21 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U7  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n16 ), .A2(
        CipherErrorVec[33]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n17 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U6  ( .A(
        AddRoundKeyOutput[44]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n15 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U5  ( .A1(
        CipherErrorVec[33]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n14 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n15 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U4  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n16 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n14 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U3  ( .A1(
        CipherErrorVec[34]), .A2(CipherErrorVec[35]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n16 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U19  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n32 ), .ZN(
        PermutationInput[46]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n29 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n30 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U15  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n25 ), .B(
        AddRoundKeyOutput[46]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n29 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U14  ( .A1(
        CipherErrorVec[34]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n24 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U13  ( .A1(
        CipherErrorVec[35]), .A2(CipherErrorVec[33]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n24 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U12  ( .A(
        AddRoundKeyOutput[45]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n23 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U11  ( .A1(
        CipherErrorVec[35]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n23 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n33 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U9  ( .A(
        AddRoundKeyOutput[44]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n21 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U7  ( .A1(
        CipherErrorVec[34]), .A2(CipherErrorVec[33]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n22 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U6  ( .A(
        CipherErrorVec[35]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n20 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U5  ( .A(
        AddRoundKeyOutput[47]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n19 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n27 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U4  ( .A1(
        CipherErrorVec[33]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U3  ( .A1(
        CipherErrorVec[35]), .A2(CipherErrorVec[34]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n18 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U26  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n48 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n47 ), .ZN(
        PermutationInput[47]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U25  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n46 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n45 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n47 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n44 ), .A2(
        AddRoundKeyOutput[44]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n45 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n43 ), .A2(
        AddRoundKeyOutput[47]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n46 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n42 ), .A2(
        CipherErrorVec[33]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n40 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n48 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U20  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n39 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n38 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n40 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U19  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n44 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n38 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n42 ), .A2(
        AddRoundKeyOutput[47]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n44 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U17  ( .A1(
        CipherErrorVec[33]), .A2(AddRoundKeyOutput[44]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n39 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n37 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n36 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U14  ( .A1(
        CipherErrorVec[33]), .A2(AddRoundKeyOutput[47]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U13  ( .A(
        AddRoundKeyOutput[46]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n33 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n35 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U12  ( .A1(
        CipherErrorVec[34]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n33 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U11  ( .A(
        CipherErrorVec[35]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n29 ), .A2(
        AddRoundKeyOutput[46]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n30 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U8  ( .A1(
        CipherErrorVec[33]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n29 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U7  ( .A(
        AddRoundKeyOutput[47]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n42 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n28 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U6  ( .A1(
        CipherErrorVec[34]), .A2(CipherErrorVec[35]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n42 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n27 ), .B(
        AddRoundKeyOutput[45]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U4  ( .A1(
        CipherErrorVec[35]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U3  ( .A1(
        CipherErrorVec[34]), .A2(CipherErrorVec[33]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n44 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n43 ), .ZN(
        PermutationInput[48]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n42 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n41 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n40 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n39 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n44 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n38 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n37 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n39 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U20  ( .A1(
        AddRoundKeyOutput[48]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U19  ( .A1(
        CipherErrorVec[38]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n35 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n36 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U18  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n38 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n40 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U16  ( .A1(
        CipherErrorVec[38]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n31 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n32 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U15  ( .A1(
        AddRoundKeyOutput[48]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n31 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n30 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n42 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U12  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n29 ), .B(
        AddRoundKeyOutput[50]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n42 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U11  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n28 ), .A2(
        CipherErrorVec[37]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n29 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U10  ( .A1(
        CipherErrorVec[38]), .A2(CipherErrorVec[36]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U9  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n27 ), .B(
        AddRoundKeyOutput[51]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n26 ), .A2(
        CipherErrorVec[36]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U7  ( .A1(
        CipherErrorVec[38]), .A2(CipherErrorVec[37]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n26 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U6  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n35 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n24 ), .B(
        AddRoundKeyOutput[49]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n33 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U4  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n25 ), .A2(
        CipherErrorVec[38]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U3  ( .A1(
        CipherErrorVec[36]), .A2(CipherErrorVec[37]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n25 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n24 ), .ZN(
        PermutationInput[49]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n23 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n21 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n20 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n22 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U12  ( .A(
        AddRoundKeyOutput[50]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n19 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n23 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U11  ( .A1(
        CipherErrorVec[37]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U10  ( .A1(
        CipherErrorVec[36]), .A2(CipherErrorVec[38]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n18 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U8  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n17 ), .B(
        AddRoundKeyOutput[51]), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n21 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U7  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n16 ), .A2(
        CipherErrorVec[36]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n17 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U6  ( .A(
        AddRoundKeyOutput[48]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n15 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U5  ( .A1(
        CipherErrorVec[36]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n14 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n15 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U4  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n16 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n14 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U3  ( .A1(
        CipherErrorVec[37]), .A2(CipherErrorVec[38]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n16 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U19  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n32 ), .ZN(
        PermutationInput[50]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n29 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n30 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U15  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n25 ), .B(
        AddRoundKeyOutput[50]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n29 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U14  ( .A1(
        CipherErrorVec[37]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n24 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U13  ( .A1(
        CipherErrorVec[38]), .A2(CipherErrorVec[36]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n24 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U12  ( .A(
        AddRoundKeyOutput[49]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n23 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U11  ( .A1(
        CipherErrorVec[38]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n23 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n33 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U9  ( .A(
        AddRoundKeyOutput[48]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n21 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U7  ( .A1(
        CipherErrorVec[37]), .A2(CipherErrorVec[36]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n22 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U6  ( .A(
        CipherErrorVec[38]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n20 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U5  ( .A(
        AddRoundKeyOutput[51]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n19 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n27 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U4  ( .A1(
        CipherErrorVec[36]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U3  ( .A1(
        CipherErrorVec[38]), .A2(CipherErrorVec[37]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n18 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U26  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n48 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n47 ), .ZN(
        PermutationInput[51]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U25  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n46 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n45 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n47 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n44 ), .A2(
        AddRoundKeyOutput[48]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n45 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n43 ), .A2(
        AddRoundKeyOutput[51]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n46 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n42 ), .A2(
        CipherErrorVec[36]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n40 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n48 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U20  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n39 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n38 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n40 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U19  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n44 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n38 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n42 ), .A2(
        AddRoundKeyOutput[51]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n44 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U17  ( .A1(
        CipherErrorVec[36]), .A2(AddRoundKeyOutput[48]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n39 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n37 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n36 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U14  ( .A1(
        CipherErrorVec[36]), .A2(AddRoundKeyOutput[51]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U13  ( .A(
        AddRoundKeyOutput[50]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n33 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n35 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U12  ( .A1(
        CipherErrorVec[37]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n33 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U11  ( .A(
        CipherErrorVec[38]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n29 ), .A2(
        AddRoundKeyOutput[50]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n30 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U8  ( .A1(
        CipherErrorVec[36]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n29 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U7  ( .A(
        AddRoundKeyOutput[51]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n42 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n28 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U6  ( .A1(
        CipherErrorVec[37]), .A2(CipherErrorVec[38]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n42 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n27 ), .B(
        AddRoundKeyOutput[49]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U4  ( .A1(
        CipherErrorVec[38]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U3  ( .A1(
        CipherErrorVec[37]), .A2(CipherErrorVec[36]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n44 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n43 ), .ZN(
        PermutationInput[52]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n42 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n41 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n40 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n39 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n44 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n38 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n37 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n39 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U20  ( .A1(
        AddRoundKeyOutput[52]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U19  ( .A1(
        CipherErrorVec[41]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n35 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n36 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U18  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n38 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n40 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U16  ( .A1(
        CipherErrorVec[41]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n31 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n32 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U15  ( .A1(
        AddRoundKeyOutput[52]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n31 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n30 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n42 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U12  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n29 ), .B(
        AddRoundKeyOutput[54]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n42 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U11  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n28 ), .A2(
        CipherErrorVec[40]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n29 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U10  ( .A1(
        CipherErrorVec[41]), .A2(CipherErrorVec[39]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U9  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n27 ), .B(
        AddRoundKeyOutput[55]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n26 ), .A2(
        CipherErrorVec[39]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U7  ( .A1(
        CipherErrorVec[41]), .A2(CipherErrorVec[40]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n26 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U6  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n35 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n24 ), .B(
        AddRoundKeyOutput[53]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n33 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U4  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n25 ), .A2(
        CipherErrorVec[41]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U3  ( .A1(
        CipherErrorVec[39]), .A2(CipherErrorVec[40]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n25 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n24 ), .ZN(
        PermutationInput[53]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n23 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n21 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n20 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n22 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U12  ( .A(
        AddRoundKeyOutput[54]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n19 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n23 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U11  ( .A1(
        CipherErrorVec[40]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U10  ( .A1(
        CipherErrorVec[39]), .A2(CipherErrorVec[41]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n18 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U8  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n17 ), .B(
        AddRoundKeyOutput[55]), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n21 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U7  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n16 ), .A2(
        CipherErrorVec[39]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n17 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U6  ( .A(
        AddRoundKeyOutput[52]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n15 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U5  ( .A1(
        CipherErrorVec[39]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n14 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n15 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U4  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n16 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n14 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U3  ( .A1(
        CipherErrorVec[40]), .A2(CipherErrorVec[41]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n16 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U19  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n32 ), .ZN(
        PermutationInput[54]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n29 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n30 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U15  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n25 ), .B(
        AddRoundKeyOutput[54]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n29 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U14  ( .A1(
        CipherErrorVec[40]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n24 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U13  ( .A1(
        CipherErrorVec[41]), .A2(CipherErrorVec[39]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n24 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U12  ( .A(
        AddRoundKeyOutput[53]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n23 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U11  ( .A1(
        CipherErrorVec[41]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n23 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n33 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U9  ( .A(
        AddRoundKeyOutput[52]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n21 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U7  ( .A1(
        CipherErrorVec[40]), .A2(CipherErrorVec[39]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n22 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U6  ( .A(
        CipherErrorVec[41]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n20 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U5  ( .A(
        AddRoundKeyOutput[55]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n19 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n27 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U4  ( .A1(
        CipherErrorVec[39]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U3  ( .A1(
        CipherErrorVec[41]), .A2(CipherErrorVec[40]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n18 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U26  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n48 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n47 ), .ZN(
        PermutationInput[55]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U25  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n46 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n45 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n47 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n44 ), .A2(
        AddRoundKeyOutput[52]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n45 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n43 ), .A2(
        AddRoundKeyOutput[55]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n46 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n42 ), .A2(
        CipherErrorVec[39]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n40 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n48 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U20  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n39 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n38 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n40 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U19  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n44 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n38 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n42 ), .A2(
        AddRoundKeyOutput[55]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n44 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U17  ( .A1(
        CipherErrorVec[39]), .A2(AddRoundKeyOutput[52]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n39 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n37 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n36 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U14  ( .A1(
        CipherErrorVec[39]), .A2(AddRoundKeyOutput[55]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U13  ( .A(
        AddRoundKeyOutput[54]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n33 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n35 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U12  ( .A1(
        CipherErrorVec[40]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n33 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U11  ( .A(
        CipherErrorVec[41]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n29 ), .A2(
        AddRoundKeyOutput[54]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n30 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U8  ( .A1(
        CipherErrorVec[39]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n29 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U7  ( .A(
        AddRoundKeyOutput[55]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n42 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n28 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U6  ( .A1(
        CipherErrorVec[40]), .A2(CipherErrorVec[41]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n42 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n27 ), .B(
        AddRoundKeyOutput[53]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U4  ( .A1(
        CipherErrorVec[41]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U3  ( .A1(
        CipherErrorVec[40]), .A2(CipherErrorVec[39]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n44 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n43 ), .ZN(
        PermutationInput[56]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n42 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n41 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n40 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n39 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n44 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n38 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n37 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n39 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U20  ( .A1(
        AddRoundKeyOutput[56]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U19  ( .A1(
        CipherErrorVec[44]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n35 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n36 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U18  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n38 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n40 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U16  ( .A1(
        CipherErrorVec[44]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n31 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n32 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U15  ( .A1(
        AddRoundKeyOutput[56]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n31 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n30 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n42 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U12  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n29 ), .B(
        AddRoundKeyOutput[58]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n42 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U11  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n28 ), .A2(
        CipherErrorVec[43]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n29 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U10  ( .A1(
        CipherErrorVec[44]), .A2(CipherErrorVec[42]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U9  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n27 ), .B(
        AddRoundKeyOutput[59]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n26 ), .A2(
        CipherErrorVec[42]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U7  ( .A1(
        CipherErrorVec[44]), .A2(CipherErrorVec[43]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n26 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U6  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n35 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n24 ), .B(
        AddRoundKeyOutput[57]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n33 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U4  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n25 ), .A2(
        CipherErrorVec[44]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U3  ( .A1(
        CipherErrorVec[42]), .A2(CipherErrorVec[43]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n25 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n24 ), .ZN(
        PermutationInput[57]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n23 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n21 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n20 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n22 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U12  ( .A(
        AddRoundKeyOutput[58]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n19 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n23 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U11  ( .A1(
        CipherErrorVec[43]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U10  ( .A1(
        CipherErrorVec[42]), .A2(CipherErrorVec[44]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n18 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U8  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n17 ), .B(
        AddRoundKeyOutput[59]), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n21 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U7  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n16 ), .A2(
        CipherErrorVec[42]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n17 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U6  ( .A(
        AddRoundKeyOutput[56]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n15 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U5  ( .A1(
        CipherErrorVec[42]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n14 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n15 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U4  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n16 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n14 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U3  ( .A1(
        CipherErrorVec[43]), .A2(CipherErrorVec[44]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n16 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U19  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n32 ), .ZN(
        PermutationInput[58]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n29 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n30 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U15  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n25 ), .B(
        AddRoundKeyOutput[58]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n29 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U14  ( .A1(
        CipherErrorVec[43]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n24 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U13  ( .A1(
        CipherErrorVec[44]), .A2(CipherErrorVec[42]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n24 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U12  ( .A(
        AddRoundKeyOutput[57]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n23 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U11  ( .A1(
        CipherErrorVec[44]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n23 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n33 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U9  ( .A(
        AddRoundKeyOutput[56]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n21 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U7  ( .A1(
        CipherErrorVec[43]), .A2(CipherErrorVec[42]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n22 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U6  ( .A(
        CipherErrorVec[44]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n20 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U5  ( .A(
        AddRoundKeyOutput[59]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n19 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n27 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U4  ( .A1(
        CipherErrorVec[42]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U3  ( .A1(
        CipherErrorVec[44]), .A2(CipherErrorVec[43]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n18 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U26  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n48 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n47 ), .ZN(
        PermutationInput[59]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U25  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n46 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n45 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n47 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n44 ), .A2(
        AddRoundKeyOutput[56]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n45 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n43 ), .A2(
        AddRoundKeyOutput[59]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n46 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n42 ), .A2(
        CipherErrorVec[42]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n40 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n48 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U20  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n39 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n38 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n40 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U19  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n44 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n38 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n42 ), .A2(
        AddRoundKeyOutput[59]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n44 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U17  ( .A1(
        CipherErrorVec[42]), .A2(AddRoundKeyOutput[56]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n39 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n37 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n36 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U14  ( .A1(
        CipherErrorVec[42]), .A2(AddRoundKeyOutput[59]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U13  ( .A(
        AddRoundKeyOutput[58]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n33 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n35 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U12  ( .A1(
        CipherErrorVec[43]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n33 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U11  ( .A(
        CipherErrorVec[44]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n29 ), .A2(
        AddRoundKeyOutput[58]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n30 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U8  ( .A1(
        CipherErrorVec[42]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n29 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U7  ( .A(
        AddRoundKeyOutput[59]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n42 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n28 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U6  ( .A1(
        CipherErrorVec[43]), .A2(CipherErrorVec[44]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n42 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n27 ), .B(
        AddRoundKeyOutput[57]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U4  ( .A1(
        CipherErrorVec[44]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U3  ( .A1(
        CipherErrorVec[43]), .A2(CipherErrorVec[42]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n44 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n43 ), .ZN(
        PermutationInput[60]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n42 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n41 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n40 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n39 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n44 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n38 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n37 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n39 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U20  ( .A1(
        AddRoundKeyOutput[60]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U19  ( .A1(
        CipherErrorVec[47]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n35 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n36 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U18  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n38 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n40 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U16  ( .A1(
        CipherErrorVec[47]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n31 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n32 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U15  ( .A1(
        AddRoundKeyOutput[60]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n31 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n30 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n42 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U12  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n29 ), .B(
        AddRoundKeyOutput[62]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n42 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U11  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n28 ), .A2(
        CipherErrorVec[46]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n29 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U10  ( .A1(
        CipherErrorVec[47]), .A2(CipherErrorVec[45]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U9  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n27 ), .B(
        AddRoundKeyOutput[63]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n26 ), .A2(
        CipherErrorVec[45]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U7  ( .A1(
        CipherErrorVec[47]), .A2(CipherErrorVec[46]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n26 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U6  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n35 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n24 ), .B(
        AddRoundKeyOutput[61]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n33 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U4  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n25 ), .A2(
        CipherErrorVec[47]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U3  ( .A1(
        CipherErrorVec[45]), .A2(CipherErrorVec[46]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n25 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n24 ), .ZN(
        PermutationInput[61]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U14  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n23 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U13  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n21 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n20 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n22 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U12  ( .A(
        AddRoundKeyOutput[62]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n19 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n23 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U11  ( .A1(
        CipherErrorVec[46]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U10  ( .A1(
        CipherErrorVec[45]), .A2(CipherErrorVec[47]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n18 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U8  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n17 ), .B(
        AddRoundKeyOutput[63]), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n21 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U7  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n16 ), .A2(
        CipherErrorVec[45]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n17 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U6  ( .A(
        AddRoundKeyOutput[60]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n15 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U5  ( .A1(
        CipherErrorVec[45]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n14 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n15 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U4  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n16 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n14 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U3  ( .A1(
        CipherErrorVec[46]), .A2(CipherErrorVec[47]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n16 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U19  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n33 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n32 ), .ZN(
        PermutationInput[62]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U17  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n29 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n30 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n28 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U15  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n25 ), .B(
        AddRoundKeyOutput[62]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n29 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U14  ( .A1(
        CipherErrorVec[46]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n24 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n25 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U13  ( .A1(
        CipherErrorVec[47]), .A2(CipherErrorVec[45]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n24 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U12  ( .A(
        AddRoundKeyOutput[61]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n23 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U11  ( .A1(
        CipherErrorVec[47]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n23 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n27 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n33 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U9  ( .A(
        AddRoundKeyOutput[60]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n26 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U8  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n20 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n22 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n21 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U7  ( .A1(
        CipherErrorVec[46]), .A2(CipherErrorVec[45]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n22 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U6  ( .A(
        CipherErrorVec[47]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n20 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U5  ( .A(
        AddRoundKeyOutput[63]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n19 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n27 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U4  ( .A1(
        CipherErrorVec[45]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n18 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n19 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U3  ( .A1(
        CipherErrorVec[47]), .A2(CipherErrorVec[46]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n18 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U26  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n48 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n47 ), .ZN(
        PermutationInput[63]) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U25  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n46 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n45 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n47 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U24  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n44 ), .A2(
        AddRoundKeyOutput[60]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n45 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U23  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n43 ), .A2(
        AddRoundKeyOutput[63]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n46 ) );
  OR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U22  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n42 ), .A2(
        CipherErrorVec[45]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n43 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U21  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n41 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n40 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n48 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U20  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n39 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n38 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n40 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U19  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n44 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n38 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U18  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n42 ), .A2(
        AddRoundKeyOutput[63]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n44 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U17  ( .A1(
        CipherErrorVec[45]), .A2(AddRoundKeyOutput[60]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n39 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U16  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n37 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n36 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n41 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U15  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n35 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n34 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n36 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U14  ( .A1(
        CipherErrorVec[45]), .A2(AddRoundKeyOutput[63]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n34 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U13  ( .A(
        AddRoundKeyOutput[62]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n33 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n35 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U12  ( .A1(
        CipherErrorVec[46]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n32 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n33 ) );
  INV_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U11  ( .A(
        CipherErrorVec[47]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n32 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U10  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n31 ), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n30 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n37 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U9  ( .A1(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n29 ), .A2(
        AddRoundKeyOutput[62]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n30 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U8  ( .A1(
        CipherErrorVec[45]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n28 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n29 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U7  ( .A(
        AddRoundKeyOutput[63]), .B(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n42 ), .Z(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n28 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U6  ( .A1(
        CipherErrorVec[46]), .A2(CipherErrorVec[47]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n42 ) );
  XNOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U5  ( .A(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n27 ), .B(
        AddRoundKeyOutput[61]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n31 ) );
  NOR2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U4  ( .A1(
        CipherErrorVec[47]), .A2(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n27 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U3  ( .A1(
        CipherErrorVec[46]), .A2(CipherErrorVec[45]), .ZN(
        \SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n26 ) );
  DFF_X1 \StateReg_s_current_state_reg[0]  ( .D(PermutationInput[0]), .CK(clk), 
        .Q(Feedback[60]) );
  DFF_X1 \StateReg_s_current_state_reg[1]  ( .D(PermutationInput[1]), .CK(clk), 
        .Q(Feedback[61]) );
  DFF_X1 \StateReg_s_current_state_reg[2]  ( .D(PermutationInput[2]), .CK(clk), 
        .Q(Feedback[62]) );
  DFF_X1 \StateReg_s_current_state_reg[3]  ( .D(PermutationInput[3]), .CK(clk), 
        .Q(Feedback[63]) );
  DFF_X1 \StateReg_s_current_state_reg[4]  ( .D(PermutationInput[4]), .CK(clk), 
        .Q(Feedback[48]) );
  DFF_X1 \StateReg_s_current_state_reg[5]  ( .D(PermutationInput[5]), .CK(clk), 
        .Q(Feedback[49]) );
  DFF_X1 \StateReg_s_current_state_reg[6]  ( .D(PermutationInput[6]), .CK(clk), 
        .Q(Feedback[50]) );
  DFF_X1 \StateReg_s_current_state_reg[7]  ( .D(PermutationInput[7]), .CK(clk), 
        .Q(Feedback[51]) );
  DFF_X1 \StateReg_s_current_state_reg[8]  ( .D(PermutationInput[8]), .CK(clk), 
        .Q(Feedback[52]) );
  DFF_X1 \StateReg_s_current_state_reg[9]  ( .D(PermutationInput[9]), .CK(clk), 
        .Q(Feedback[53]) );
  DFF_X1 \StateReg_s_current_state_reg[10]  ( .D(PermutationInput[10]), .CK(
        clk), .Q(Feedback[54]) );
  DFF_X1 \StateReg_s_current_state_reg[11]  ( .D(PermutationInput[11]), .CK(
        clk), .Q(Feedback[55]) );
  DFF_X1 \StateReg_s_current_state_reg[12]  ( .D(PermutationInput[12]), .CK(
        clk), .Q(Feedback[56]) );
  DFF_X1 \StateReg_s_current_state_reg[13]  ( .D(PermutationInput[13]), .CK(
        clk), .Q(Feedback[57]) );
  DFF_X1 \StateReg_s_current_state_reg[14]  ( .D(PermutationInput[14]), .CK(
        clk), .Q(Feedback[58]) );
  DFF_X1 \StateReg_s_current_state_reg[15]  ( .D(PermutationInput[15]), .CK(
        clk), .Q(Feedback[59]) );
  DFF_X1 \StateReg_s_current_state_reg[16]  ( .D(PermutationInput[16]), .CK(
        clk), .Q(Feedback[32]) );
  DFF_X1 \StateReg_s_current_state_reg[17]  ( .D(PermutationInput[17]), .CK(
        clk), .Q(Feedback[33]) );
  DFF_X1 \StateReg_s_current_state_reg[18]  ( .D(PermutationInput[18]), .CK(
        clk), .Q(Feedback[34]) );
  DFF_X1 \StateReg_s_current_state_reg[19]  ( .D(PermutationInput[19]), .CK(
        clk), .Q(Feedback[35]) );
  DFF_X1 \StateReg_s_current_state_reg[20]  ( .D(PermutationInput[20]), .CK(
        clk), .Q(Feedback[44]) );
  DFF_X1 \StateReg_s_current_state_reg[21]  ( .D(PermutationInput[21]), .CK(
        clk), .Q(Feedback[45]) );
  DFF_X1 \StateReg_s_current_state_reg[22]  ( .D(PermutationInput[22]), .CK(
        clk), .Q(Feedback[46]) );
  DFF_X1 \StateReg_s_current_state_reg[23]  ( .D(PermutationInput[23]), .CK(
        clk), .Q(Feedback[47]) );
  DFF_X1 \StateReg_s_current_state_reg[24]  ( .D(PermutationInput[24]), .CK(
        clk), .Q(Feedback[40]) );
  DFF_X1 \StateReg_s_current_state_reg[25]  ( .D(PermutationInput[25]), .CK(
        clk), .Q(Feedback[41]) );
  DFF_X1 \StateReg_s_current_state_reg[26]  ( .D(PermutationInput[26]), .CK(
        clk), .Q(Feedback[42]) );
  DFF_X1 \StateReg_s_current_state_reg[27]  ( .D(PermutationInput[27]), .CK(
        clk), .Q(Feedback[43]) );
  DFF_X1 \StateReg_s_current_state_reg[28]  ( .D(PermutationInput[28]), .CK(
        clk), .Q(Feedback[36]) );
  DFF_X1 \StateReg_s_current_state_reg[29]  ( .D(PermutationInput[29]), .CK(
        clk), .Q(Feedback[37]) );
  DFF_X1 \StateReg_s_current_state_reg[30]  ( .D(PermutationInput[30]), .CK(
        clk), .Q(Feedback[38]) );
  DFF_X1 \StateReg_s_current_state_reg[31]  ( .D(PermutationInput[31]), .CK(
        clk), .Q(Feedback[39]) );
  DFF_X1 \StateReg_s_current_state_reg[32]  ( .D(PermutationInput[32]), .CK(
        clk), .Q(Feedback[16]) );
  DFF_X1 \StateReg_s_current_state_reg[33]  ( .D(PermutationInput[33]), .CK(
        clk), .Q(Feedback[17]) );
  DFF_X1 \StateReg_s_current_state_reg[34]  ( .D(PermutationInput[34]), .CK(
        clk), .Q(Feedback[18]) );
  DFF_X1 \StateReg_s_current_state_reg[35]  ( .D(PermutationInput[35]), .CK(
        clk), .Q(Feedback[19]) );
  DFF_X1 \StateReg_s_current_state_reg[36]  ( .D(PermutationInput[36]), .CK(
        clk), .Q(Feedback[28]) );
  DFF_X1 \StateReg_s_current_state_reg[37]  ( .D(PermutationInput[37]), .CK(
        clk), .Q(Feedback[29]) );
  DFF_X1 \StateReg_s_current_state_reg[38]  ( .D(PermutationInput[38]), .CK(
        clk), .Q(Feedback[30]) );
  DFF_X1 \StateReg_s_current_state_reg[39]  ( .D(PermutationInput[39]), .CK(
        clk), .Q(Feedback[31]) );
  DFF_X1 \StateReg_s_current_state_reg[40]  ( .D(PermutationInput[40]), .CK(
        clk), .Q(Feedback[24]) );
  DFF_X1 \StateReg_s_current_state_reg[41]  ( .D(PermutationInput[41]), .CK(
        clk), .Q(Feedback[25]) );
  DFF_X1 \StateReg_s_current_state_reg[42]  ( .D(PermutationInput[42]), .CK(
        clk), .Q(Feedback[26]) );
  DFF_X1 \StateReg_s_current_state_reg[43]  ( .D(PermutationInput[43]), .CK(
        clk), .Q(Feedback[27]) );
  DFF_X1 \StateReg_s_current_state_reg[44]  ( .D(PermutationInput[44]), .CK(
        clk), .Q(Feedback[20]) );
  DFF_X1 \StateReg_s_current_state_reg[45]  ( .D(PermutationInput[45]), .CK(
        clk), .Q(Feedback[21]) );
  DFF_X1 \StateReg_s_current_state_reg[46]  ( .D(PermutationInput[46]), .CK(
        clk), .Q(Feedback[22]) );
  DFF_X1 \StateReg_s_current_state_reg[47]  ( .D(PermutationInput[47]), .CK(
        clk), .Q(Feedback[23]) );
  DFF_X1 \StateReg_s_current_state_reg[48]  ( .D(PermutationInput[48]), .CK(
        clk), .Q(Feedback[4]) );
  DFF_X1 \StateReg_s_current_state_reg[49]  ( .D(PermutationInput[49]), .CK(
        clk), .Q(Feedback[5]) );
  DFF_X1 \StateReg_s_current_state_reg[50]  ( .D(PermutationInput[50]), .CK(
        clk), .Q(Feedback[6]) );
  DFF_X1 \StateReg_s_current_state_reg[51]  ( .D(PermutationInput[51]), .CK(
        clk), .Q(Feedback[7]) );
  DFF_X1 \StateReg_s_current_state_reg[52]  ( .D(PermutationInput[52]), .CK(
        clk), .Q(Feedback[8]) );
  DFF_X1 \StateReg_s_current_state_reg[53]  ( .D(PermutationInput[53]), .CK(
        clk), .Q(Feedback[9]) );
  DFF_X1 \StateReg_s_current_state_reg[54]  ( .D(PermutationInput[54]), .CK(
        clk), .Q(Feedback[10]) );
  DFF_X1 \StateReg_s_current_state_reg[55]  ( .D(PermutationInput[55]), .CK(
        clk), .Q(Feedback[11]) );
  DFF_X1 \StateReg_s_current_state_reg[56]  ( .D(PermutationInput[56]), .CK(
        clk), .Q(Feedback[12]) );
  DFF_X1 \StateReg_s_current_state_reg[57]  ( .D(PermutationInput[57]), .CK(
        clk), .Q(Feedback[13]) );
  DFF_X1 \StateReg_s_current_state_reg[58]  ( .D(PermutationInput[58]), .CK(
        clk), .Q(Feedback[14]) );
  DFF_X1 \StateReg_s_current_state_reg[59]  ( .D(PermutationInput[59]), .CK(
        clk), .Q(Feedback[15]) );
  DFF_X1 \StateReg_s_current_state_reg[60]  ( .D(PermutationInput[60]), .CK(
        clk), .Q(Feedback[0]) );
  DFF_X1 \StateReg_s_current_state_reg[61]  ( .D(PermutationInput[61]), .CK(
        clk), .Q(Feedback[1]) );
  DFF_X1 \StateReg_s_current_state_reg[62]  ( .D(PermutationInput[62]), .CK(
        clk), .Q(Feedback[2]) );
  DFF_X1 \StateReg_s_current_state_reg[63]  ( .D(PermutationInput[63]), .CK(
        clk), .Q(Feedback[3]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_0_LFInst_0_n2 ), .B(Input[1]), .ZN(
        Red_MCOutput[0]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_0_U3  ( .A(Input[2]), .B(
        Input[0]), .ZN(\Red_PlaintextInst_LFInst_0_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_0_LFInst_1_n2 ), .B(Input[1]), .ZN(
        Red_MCOutput[1]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_1_U3  ( .A(Input[3]), .B(
        Input[0]), .ZN(\Red_PlaintextInst_LFInst_0_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_0_LFInst_2_n2 ), .B(Input[2]), .ZN(
        Red_MCOutput[2]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_2_U3  ( .A(Input[3]), .B(
        Input[0]), .ZN(\Red_PlaintextInst_LFInst_0_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_1_LFInst_0_n2 ), .B(Input[5]), .ZN(
        Red_MCOutput[3]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_0_U3  ( .A(Input[6]), .B(
        Input[4]), .ZN(\Red_PlaintextInst_LFInst_1_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_1_LFInst_1_n2 ), .B(Input[5]), .ZN(
        Red_MCOutput[4]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_1_U3  ( .A(Input[7]), .B(
        Input[4]), .ZN(\Red_PlaintextInst_LFInst_1_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_1_LFInst_2_n2 ), .B(Input[6]), .ZN(
        Red_MCOutput[5]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_2_U3  ( .A(Input[7]), .B(
        Input[4]), .ZN(\Red_PlaintextInst_LFInst_1_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_2_LFInst_0_n2 ), .B(Input[9]), .ZN(
        Red_MCOutput[6]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_0_U3  ( .A(Input[10]), .B(
        Input[8]), .ZN(\Red_PlaintextInst_LFInst_2_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_2_LFInst_1_n2 ), .B(Input[9]), .ZN(
        Red_MCOutput[7]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_1_U3  ( .A(Input[11]), .B(
        Input[8]), .ZN(\Red_PlaintextInst_LFInst_2_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_2_LFInst_2_n2 ), .B(Input[10]), .ZN(
        Red_MCOutput[8]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_2_U3  ( .A(Input[11]), .B(
        Input[8]), .ZN(\Red_PlaintextInst_LFInst_2_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_3_LFInst_0_n2 ), .B(Input[13]), .ZN(
        Red_MCOutput[9]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_0_U3  ( .A(Input[14]), .B(
        Input[12]), .ZN(\Red_PlaintextInst_LFInst_3_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_3_LFInst_1_n2 ), .B(Input[13]), .ZN(
        Red_MCOutput[10]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_1_U3  ( .A(Input[15]), .B(
        Input[12]), .ZN(\Red_PlaintextInst_LFInst_3_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_3_LFInst_2_n2 ), .B(Input[14]), .ZN(
        Red_MCOutput[11]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_2_U3  ( .A(Input[15]), .B(
        Input[12]), .ZN(\Red_PlaintextInst_LFInst_3_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_4_LFInst_0_n2 ), .B(Input[17]), .ZN(
        Red_MCOutput[12]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_0_U3  ( .A(Input[18]), .B(
        Input[16]), .ZN(\Red_PlaintextInst_LFInst_4_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_4_LFInst_1_n2 ), .B(Input[17]), .ZN(
        Red_MCOutput[13]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_1_U3  ( .A(Input[19]), .B(
        Input[16]), .ZN(\Red_PlaintextInst_LFInst_4_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_4_LFInst_2_n2 ), .B(Input[18]), .ZN(
        Red_MCOutput[14]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_2_U3  ( .A(Input[19]), .B(
        Input[16]), .ZN(\Red_PlaintextInst_LFInst_4_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_5_LFInst_0_n2 ), .B(Input[21]), .ZN(
        Red_MCOutput[15]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_0_U3  ( .A(Input[22]), .B(
        Input[20]), .ZN(\Red_PlaintextInst_LFInst_5_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_5_LFInst_1_n2 ), .B(Input[21]), .ZN(
        Red_MCOutput[16]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_1_U3  ( .A(Input[23]), .B(
        Input[20]), .ZN(\Red_PlaintextInst_LFInst_5_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_5_LFInst_2_n2 ), .B(Input[22]), .ZN(
        Red_MCOutput[17]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_2_U3  ( .A(Input[23]), .B(
        Input[20]), .ZN(\Red_PlaintextInst_LFInst_5_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_6_LFInst_0_n2 ), .B(Input[25]), .ZN(
        Red_MCOutput[18]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_0_U3  ( .A(Input[26]), .B(
        Input[24]), .ZN(\Red_PlaintextInst_LFInst_6_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_6_LFInst_1_n2 ), .B(Input[25]), .ZN(
        Red_MCOutput[19]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_1_U3  ( .A(Input[27]), .B(
        Input[24]), .ZN(\Red_PlaintextInst_LFInst_6_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_6_LFInst_2_n2 ), .B(Input[26]), .ZN(
        Red_MCOutput[20]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_2_U3  ( .A(Input[27]), .B(
        Input[24]), .ZN(\Red_PlaintextInst_LFInst_6_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_7_LFInst_0_n2 ), .B(Input[29]), .ZN(
        Red_MCOutput[21]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_0_U3  ( .A(Input[30]), .B(
        Input[28]), .ZN(\Red_PlaintextInst_LFInst_7_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_7_LFInst_1_n2 ), .B(Input[29]), .ZN(
        Red_MCOutput[22]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_1_U3  ( .A(Input[31]), .B(
        Input[28]), .ZN(\Red_PlaintextInst_LFInst_7_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_7_LFInst_2_n2 ), .B(Input[30]), .ZN(
        Red_MCOutput[23]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_2_U3  ( .A(Input[31]), .B(
        Input[28]), .ZN(\Red_PlaintextInst_LFInst_7_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_8_LFInst_0_n2 ), .B(Input[33]), .ZN(
        Red_Input[24]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_0_U3  ( .A(Input[34]), .B(
        Input[32]), .ZN(\Red_PlaintextInst_LFInst_8_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_8_LFInst_1_n2 ), .B(Input[33]), .ZN(
        Red_Input[25]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_1_U3  ( .A(Input[35]), .B(
        Input[32]), .ZN(\Red_PlaintextInst_LFInst_8_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_8_LFInst_2_n2 ), .B(Input[34]), .ZN(
        Red_Input[26]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_2_U3  ( .A(Input[35]), .B(
        Input[32]), .ZN(\Red_PlaintextInst_LFInst_8_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_9_LFInst_0_n2 ), .B(Input[37]), .ZN(
        Red_Input[27]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_0_U3  ( .A(Input[38]), .B(
        Input[36]), .ZN(\Red_PlaintextInst_LFInst_9_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_9_LFInst_1_n2 ), .B(Input[37]), .ZN(
        Red_Input[28]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_1_U3  ( .A(Input[39]), .B(
        Input[36]), .ZN(\Red_PlaintextInst_LFInst_9_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_9_LFInst_2_n2 ), .B(Input[38]), .ZN(
        Red_Input[29]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_2_U3  ( .A(Input[39]), .B(
        Input[36]), .ZN(\Red_PlaintextInst_LFInst_9_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_10_LFInst_0_n2 ), .B(Input[41]), .ZN(
        Red_Input[30]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_0_U3  ( .A(Input[42]), .B(
        Input[40]), .ZN(\Red_PlaintextInst_LFInst_10_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_10_LFInst_1_n2 ), .B(Input[41]), .ZN(
        Red_Input[31]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_1_U3  ( .A(Input[43]), .B(
        Input[40]), .ZN(\Red_PlaintextInst_LFInst_10_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_10_LFInst_2_n2 ), .B(Input[42]), .ZN(
        Red_Input[32]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_2_U3  ( .A(Input[43]), .B(
        Input[40]), .ZN(\Red_PlaintextInst_LFInst_10_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_11_LFInst_0_n2 ), .B(Input[45]), .ZN(
        Red_Input[33]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_0_U3  ( .A(Input[46]), .B(
        Input[44]), .ZN(\Red_PlaintextInst_LFInst_11_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_11_LFInst_1_n2 ), .B(Input[45]), .ZN(
        Red_Input[34]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_1_U3  ( .A(Input[47]), .B(
        Input[44]), .ZN(\Red_PlaintextInst_LFInst_11_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_11_LFInst_2_n2 ), .B(Input[46]), .ZN(
        Red_Input[35]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_2_U3  ( .A(Input[47]), .B(
        Input[44]), .ZN(\Red_PlaintextInst_LFInst_11_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_12_LFInst_0_n2 ), .B(Input[49]), .ZN(
        Red_Input[36]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_0_U3  ( .A(Input[50]), .B(
        Input[48]), .ZN(\Red_PlaintextInst_LFInst_12_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_12_LFInst_1_n2 ), .B(Input[49]), .ZN(
        Red_Input[37]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_1_U3  ( .A(Input[51]), .B(
        Input[48]), .ZN(\Red_PlaintextInst_LFInst_12_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_12_LFInst_2_n2 ), .B(Input[50]), .ZN(
        Red_Input[38]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_2_U3  ( .A(Input[51]), .B(
        Input[48]), .ZN(\Red_PlaintextInst_LFInst_12_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_13_LFInst_0_n2 ), .B(Input[53]), .ZN(
        Red_Input[39]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_0_U3  ( .A(Input[54]), .B(
        Input[52]), .ZN(\Red_PlaintextInst_LFInst_13_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_13_LFInst_1_n2 ), .B(Input[53]), .ZN(
        Red_Input[40]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_1_U3  ( .A(Input[55]), .B(
        Input[52]), .ZN(\Red_PlaintextInst_LFInst_13_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_13_LFInst_2_n2 ), .B(Input[54]), .ZN(
        Red_Input[41]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_2_U3  ( .A(Input[55]), .B(
        Input[52]), .ZN(\Red_PlaintextInst_LFInst_13_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_14_LFInst_0_n2 ), .B(Input[57]), .ZN(
        Red_Input[42]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_0_U3  ( .A(Input[58]), .B(
        Input[56]), .ZN(\Red_PlaintextInst_LFInst_14_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_14_LFInst_1_n2 ), .B(Input[57]), .ZN(
        Red_Input[43]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_1_U3  ( .A(Input[59]), .B(
        Input[56]), .ZN(\Red_PlaintextInst_LFInst_14_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_14_LFInst_2_n2 ), .B(Input[58]), .ZN(
        Red_Input[44]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_2_U3  ( .A(Input[59]), .B(
        Input[56]), .ZN(\Red_PlaintextInst_LFInst_14_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_15_LFInst_0_n2 ), .B(Input[61]), .ZN(
        Red_Input[45]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_0_U3  ( .A(Input[62]), .B(
        Input[60]), .ZN(\Red_PlaintextInst_LFInst_15_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_15_LFInst_1_n2 ), .B(Input[61]), .ZN(
        Red_Input[46]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_1_U3  ( .A(Input[63]), .B(
        Input[60]), .ZN(\Red_PlaintextInst_LFInst_15_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_15_LFInst_2_n2 ), .B(Input[62]), .ZN(
        Red_Input[47]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_2_U3  ( .A(Input[63]), .B(
        Input[60]), .ZN(\Red_PlaintextInst_LFInst_15_LFInst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_0_U2  ( .A(\Red_MCInst_XOR_r0_Inst_0_n3 ), 
        .B(Red_MCOutput[0]), .ZN(Red_MCOutput[36]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_0_U1  ( .A(Red_Input[36]), .B(
        Red_MCOutput[12]), .ZN(\Red_MCInst_XOR_r0_Inst_0_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_0_U1  ( .A(Red_Input[24]), .B(
        Red_MCOutput[0]), .Z(Red_MCOutput[24]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_1_U2  ( .A(\Red_MCInst_XOR_r0_Inst_1_n3 ), 
        .B(Red_MCOutput[1]), .ZN(Red_MCOutput[37]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_1_U1  ( .A(Red_Input[37]), .B(
        Red_MCOutput[13]), .ZN(\Red_MCInst_XOR_r0_Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_1_U1  ( .A(Red_Input[25]), .B(
        Red_MCOutput[1]), .Z(Red_MCOutput[25]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_2_U2  ( .A(\Red_MCInst_XOR_r0_Inst_2_n3 ), 
        .B(Red_MCOutput[2]), .ZN(Red_MCOutput[38]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_2_U1  ( .A(Red_Input[38]), .B(
        Red_MCOutput[14]), .ZN(\Red_MCInst_XOR_r0_Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_2_U1  ( .A(Red_Input[26]), .B(
        Red_MCOutput[2]), .Z(Red_MCOutput[26]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_3_U2  ( .A(\Red_MCInst_XOR_r0_Inst_3_n3 ), 
        .B(Red_MCOutput[3]), .ZN(Red_MCOutput[39]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_3_U1  ( .A(Red_Input[39]), .B(
        Red_MCOutput[15]), .ZN(\Red_MCInst_XOR_r0_Inst_3_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_3_U1  ( .A(Red_Input[27]), .B(
        Red_MCOutput[3]), .Z(Red_MCOutput[27]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_4_U2  ( .A(\Red_MCInst_XOR_r0_Inst_4_n3 ), 
        .B(Red_MCOutput[4]), .ZN(Red_MCOutput[40]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_4_U1  ( .A(Red_Input[40]), .B(
        Red_MCOutput[16]), .ZN(\Red_MCInst_XOR_r0_Inst_4_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_4_U1  ( .A(Red_Input[28]), .B(
        Red_MCOutput[4]), .Z(Red_MCOutput[28]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_5_U2  ( .A(\Red_MCInst_XOR_r0_Inst_5_n3 ), 
        .B(Red_MCOutput[5]), .ZN(Red_MCOutput[41]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_5_U1  ( .A(Red_Input[41]), .B(
        Red_MCOutput[17]), .ZN(\Red_MCInst_XOR_r0_Inst_5_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_5_U1  ( .A(Red_Input[29]), .B(
        Red_MCOutput[5]), .Z(Red_MCOutput[29]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_6_U2  ( .A(\Red_MCInst_XOR_r0_Inst_6_n3 ), 
        .B(Red_MCOutput[6]), .ZN(Red_MCOutput[42]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_6_U1  ( .A(Red_Input[42]), .B(
        Red_MCOutput[18]), .ZN(\Red_MCInst_XOR_r0_Inst_6_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_6_U1  ( .A(Red_Input[30]), .B(
        Red_MCOutput[6]), .Z(Red_MCOutput[30]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_7_U2  ( .A(\Red_MCInst_XOR_r0_Inst_7_n3 ), 
        .B(Red_MCOutput[7]), .ZN(Red_MCOutput[43]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_7_U1  ( .A(Red_Input[43]), .B(
        Red_MCOutput[19]), .ZN(\Red_MCInst_XOR_r0_Inst_7_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_7_U1  ( .A(Red_Input[31]), .B(
        Red_MCOutput[7]), .Z(Red_MCOutput[31]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_8_U2  ( .A(\Red_MCInst_XOR_r0_Inst_8_n3 ), 
        .B(Red_MCOutput[8]), .ZN(Red_MCOutput[44]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_8_U1  ( .A(Red_Input[44]), .B(
        Red_MCOutput[20]), .ZN(\Red_MCInst_XOR_r0_Inst_8_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_8_U1  ( .A(Red_Input[32]), .B(
        Red_MCOutput[8]), .Z(Red_MCOutput[32]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_9_U2  ( .A(\Red_MCInst_XOR_r0_Inst_9_n3 ), 
        .B(Red_MCOutput[9]), .ZN(Red_MCOutput[45]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_9_U1  ( .A(Red_Input[45]), .B(
        Red_MCOutput[21]), .ZN(\Red_MCInst_XOR_r0_Inst_9_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_9_U1  ( .A(Red_Input[33]), .B(
        Red_MCOutput[9]), .Z(Red_MCOutput[33]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_10_U2  ( .A(\Red_MCInst_XOR_r0_Inst_10_n3 ), 
        .B(Red_MCOutput[10]), .ZN(Red_MCOutput[46]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_10_U1  ( .A(Red_Input[46]), .B(
        Red_MCOutput[22]), .ZN(\Red_MCInst_XOR_r0_Inst_10_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_10_U1  ( .A(Red_Input[34]), .B(
        Red_MCOutput[10]), .Z(Red_MCOutput[34]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_11_U2  ( .A(\Red_MCInst_XOR_r0_Inst_11_n3 ), 
        .B(Red_MCOutput[11]), .ZN(Red_MCOutput[47]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_11_U1  ( .A(Red_Input[47]), .B(
        Red_MCOutput[23]), .ZN(\Red_MCInst_XOR_r0_Inst_11_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_11_U1  ( .A(Red_Input[35]), .B(
        Red_MCOutput[11]), .Z(Red_MCOutput[35]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_0_0_U1  ( .A(Red_MCOutput[36]), .B(
        Red_K0[36]), .Z(Red_AddRoundKeyOutput[36]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_0_1_U1  ( .A(Red_MCOutput[37]), .B(
        Red_K0[37]), .Z(Red_AddRoundKeyOutput[37]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_0_2_U1  ( .A(Red_MCOutput[38]), .B(
        Red_K0[38]), .Z(Red_AddRoundKeyOutput[38]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_1_0_U1  ( .A(Red_MCOutput[39]), .B(
        Red_K0[39]), .Z(Red_AddRoundKeyOutput[39]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_1_1_U1  ( .A(Red_MCOutput[40]), .B(
        Red_K0[40]), .Z(Red_AddRoundKeyOutput[40]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_1_2_U1  ( .A(Red_MCOutput[41]), .B(
        Red_K0[41]), .Z(Red_AddRoundKeyOutput[41]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_2_0_U1  ( .A(Red_MCOutput[42]), .B(
        Red_K0[42]), .Z(Red_AddRoundKeyOutput[42]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_2_1_U1  ( .A(Red_MCOutput[43]), .B(
        Red_K0[43]), .Z(Red_AddRoundKeyOutput[43]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_2_2_U1  ( .A(Red_MCOutput[44]), .B(
        Red_K0[44]), .Z(Red_AddRoundKeyOutput[44]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_3_0_U1  ( .A(Red_MCOutput[45]), .B(
        Red_K0[45]), .Z(Red_AddRoundKeyOutput[45]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_3_1_U1  ( .A(Red_MCOutput[46]), .B(
        Red_K0[46]), .Z(Red_AddRoundKeyOutput[46]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_3_2_U1  ( .A(Red_MCOutput[47]), .B(
        Red_K0[47]), .Z(Red_AddRoundKeyOutput[47]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_0_0_U1  ( .A(Red_K0[30]), .B(
        Red_MCOutput[30]), .Z(Red_AddRoundKeyOutput[30]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_0_1_U1  ( .A(Red_K0[31]), .B(
        Red_MCOutput[31]), .Z(Red_AddRoundKeyOutput[31]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_0_2_U1  ( .A(Red_K0[32]), .B(
        Red_MCOutput[32]), .Z(Red_AddRoundKeyOutput[32]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_1_0_U1  ( .A(Red_K0[33]), .B(
        Red_MCOutput[33]), .Z(Red_AddRoundKeyOutput[33]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_1_1_U1  ( .A(Red_K0[34]), .B(
        Red_MCOutput[34]), .Z(Red_AddRoundKeyOutput[34]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_1_2_U1  ( .A(Red_K0[35]), .B(
        Red_MCOutput[35]), .Z(Red_AddRoundKeyOutput[35]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_0_0_U1  ( .A(Red_MCOutput[0]), .B(Red_K0[0]), 
        .Z(Red_AddRoundKeyOutput[0]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_0_1_U1  ( .A(Red_MCOutput[1]), .B(Red_K0[1]), 
        .Z(Red_AddRoundKeyOutput[1]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_0_2_U1  ( .A(Red_MCOutput[2]), .B(Red_K0[2]), 
        .Z(Red_AddRoundKeyOutput[2]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_1_0_U1  ( .A(Red_MCOutput[3]), .B(Red_K0[3]), 
        .Z(Red_AddRoundKeyOutput[3]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_1_1_U1  ( .A(Red_MCOutput[4]), .B(Red_K0[4]), 
        .Z(Red_AddRoundKeyOutput[4]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_1_2_U1  ( .A(Red_MCOutput[5]), .B(Red_K0[5]), 
        .Z(Red_AddRoundKeyOutput[5]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_2_0_U1  ( .A(Red_MCOutput[6]), .B(Red_K0[6]), 
        .Z(Red_AddRoundKeyOutput[6]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_2_1_U1  ( .A(Red_MCOutput[7]), .B(Red_K0[7]), 
        .Z(Red_AddRoundKeyOutput[7]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_2_2_U1  ( .A(Red_MCOutput[8]), .B(Red_K0[8]), 
        .Z(Red_AddRoundKeyOutput[8]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_3_0_U1  ( .A(Red_MCOutput[9]), .B(Red_K0[9]), 
        .Z(Red_AddRoundKeyOutput[9]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_3_1_U1  ( .A(Red_MCOutput[10]), .B(
        Red_K0[10]), .Z(Red_AddRoundKeyOutput[10]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_3_2_U1  ( .A(Red_MCOutput[11]), .B(
        Red_K0[11]), .Z(Red_AddRoundKeyOutput[11]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_4_0_U1  ( .A(Red_MCOutput[12]), .B(
        Red_K0[12]), .Z(Red_AddRoundKeyOutput[12]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_4_1_U1  ( .A(Red_MCOutput[13]), .B(
        Red_K0[13]), .Z(Red_AddRoundKeyOutput[13]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_4_2_U1  ( .A(Red_MCOutput[14]), .B(
        Red_K0[14]), .Z(Red_AddRoundKeyOutput[14]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_5_0_U1  ( .A(Red_MCOutput[15]), .B(
        Red_K0[15]), .Z(Red_AddRoundKeyOutput[15]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_5_1_U1  ( .A(Red_MCOutput[16]), .B(
        Red_K0[16]), .Z(Red_AddRoundKeyOutput[16]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_5_2_U1  ( .A(Red_MCOutput[17]), .B(
        Red_K0[17]), .Z(Red_AddRoundKeyOutput[17]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_6_0_U1  ( .A(Red_MCOutput[18]), .B(
        Red_K0[18]), .Z(Red_AddRoundKeyOutput[18]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_6_1_U1  ( .A(Red_MCOutput[19]), .B(
        Red_K0[19]), .Z(Red_AddRoundKeyOutput[19]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_6_2_U1  ( .A(Red_MCOutput[20]), .B(
        Red_K0[20]), .Z(Red_AddRoundKeyOutput[20]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_7_0_U1  ( .A(Red_MCOutput[21]), .B(
        Red_K0[21]), .Z(Red_AddRoundKeyOutput[21]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_7_1_U1  ( .A(Red_MCOutput[22]), .B(
        Red_K0[22]), .Z(Red_AddRoundKeyOutput[22]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_7_2_U1  ( .A(Red_MCOutput[23]), .B(
        Red_K0[23]), .Z(Red_AddRoundKeyOutput[23]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_8_0_U1  ( .A(Red_MCOutput[24]), .B(
        Red_K0[24]), .Z(Red_AddRoundKeyOutput[24]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_8_1_U1  ( .A(Red_MCOutput[25]), .B(
        Red_K0[25]), .Z(Red_AddRoundKeyOutput[25]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_8_2_U1  ( .A(Red_MCOutput[26]), .B(
        Red_K0[26]), .Z(Red_AddRoundKeyOutput[26]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_9_0_U1  ( .A(Red_MCOutput[27]), .B(
        Red_K0[27]), .Z(Red_AddRoundKeyOutput[27]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_9_1_U1  ( .A(Red_MCOutput[28]), .B(
        Red_K0[28]), .Z(Red_AddRoundKeyOutput[28]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_9_2_U1  ( .A(Red_MCOutput[29]), .B(
        Red_K0[29]), .Z(Red_AddRoundKeyOutput[29]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_0_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst_LFInst_0_LFInst_0_n2 ), .B(AddRoundKeyOutput[1]), 
        .ZN(StateRegOutputF[0]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_0_LFInst_0_U3  ( .A(
        AddRoundKeyOutput[2]), .B(AddRoundKeyOutput[0]), .ZN(
        \StateRegOutputF_inst_LFInst_0_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_0_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst_LFInst_0_LFInst_1_n2 ), .B(AddRoundKeyOutput[1]), 
        .ZN(StateRegOutputF[1]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_0_LFInst_1_U3  ( .A(
        AddRoundKeyOutput[3]), .B(AddRoundKeyOutput[0]), .ZN(
        \StateRegOutputF_inst_LFInst_0_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_0_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst_LFInst_0_LFInst_2_n2 ), .B(AddRoundKeyOutput[2]), 
        .ZN(StateRegOutputF[2]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_0_LFInst_2_U3  ( .A(
        AddRoundKeyOutput[3]), .B(AddRoundKeyOutput[0]), .ZN(
        \StateRegOutputF_inst_LFInst_0_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_1_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst_LFInst_1_LFInst_0_n2 ), .B(AddRoundKeyOutput[5]), 
        .ZN(StateRegOutputF[3]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_1_LFInst_0_U3  ( .A(
        AddRoundKeyOutput[6]), .B(AddRoundKeyOutput[4]), .ZN(
        \StateRegOutputF_inst_LFInst_1_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_1_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst_LFInst_1_LFInst_1_n2 ), .B(AddRoundKeyOutput[5]), 
        .ZN(StateRegOutputF[4]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_1_LFInst_1_U3  ( .A(
        AddRoundKeyOutput[7]), .B(AddRoundKeyOutput[4]), .ZN(
        \StateRegOutputF_inst_LFInst_1_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_1_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst_LFInst_1_LFInst_2_n2 ), .B(AddRoundKeyOutput[6]), 
        .ZN(StateRegOutputF[5]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_1_LFInst_2_U3  ( .A(
        AddRoundKeyOutput[7]), .B(AddRoundKeyOutput[4]), .ZN(
        \StateRegOutputF_inst_LFInst_1_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_2_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst_LFInst_2_LFInst_0_n2 ), .B(AddRoundKeyOutput[9]), 
        .ZN(StateRegOutputF[6]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_2_LFInst_0_U3  ( .A(
        AddRoundKeyOutput[10]), .B(AddRoundKeyOutput[8]), .ZN(
        \StateRegOutputF_inst_LFInst_2_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_2_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst_LFInst_2_LFInst_1_n2 ), .B(AddRoundKeyOutput[9]), 
        .ZN(StateRegOutputF[7]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_2_LFInst_1_U3  ( .A(
        AddRoundKeyOutput[11]), .B(AddRoundKeyOutput[8]), .ZN(
        \StateRegOutputF_inst_LFInst_2_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_2_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst_LFInst_2_LFInst_2_n2 ), .B(AddRoundKeyOutput[10]), .ZN(StateRegOutputF[8]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_2_LFInst_2_U3  ( .A(
        AddRoundKeyOutput[11]), .B(AddRoundKeyOutput[8]), .ZN(
        \StateRegOutputF_inst_LFInst_2_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_3_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst_LFInst_3_LFInst_0_n2 ), .B(AddRoundKeyOutput[13]), .ZN(StateRegOutputF[9]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_3_LFInst_0_U3  ( .A(
        AddRoundKeyOutput[14]), .B(AddRoundKeyOutput[12]), .ZN(
        \StateRegOutputF_inst_LFInst_3_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_3_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst_LFInst_3_LFInst_1_n2 ), .B(AddRoundKeyOutput[13]), .ZN(StateRegOutputF[10]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_3_LFInst_1_U3  ( .A(
        AddRoundKeyOutput[15]), .B(AddRoundKeyOutput[12]), .ZN(
        \StateRegOutputF_inst_LFInst_3_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_3_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst_LFInst_3_LFInst_2_n2 ), .B(AddRoundKeyOutput[14]), .ZN(StateRegOutputF[11]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_3_LFInst_2_U3  ( .A(
        AddRoundKeyOutput[15]), .B(AddRoundKeyOutput[12]), .ZN(
        \StateRegOutputF_inst_LFInst_3_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_4_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst_LFInst_4_LFInst_0_n2 ), .B(AddRoundKeyOutput[17]), .ZN(StateRegOutputF[12]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_4_LFInst_0_U3  ( .A(
        AddRoundKeyOutput[18]), .B(AddRoundKeyOutput[16]), .ZN(
        \StateRegOutputF_inst_LFInst_4_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_4_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst_LFInst_4_LFInst_1_n2 ), .B(AddRoundKeyOutput[17]), .ZN(StateRegOutputF[13]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_4_LFInst_1_U3  ( .A(
        AddRoundKeyOutput[19]), .B(AddRoundKeyOutput[16]), .ZN(
        \StateRegOutputF_inst_LFInst_4_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_4_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst_LFInst_4_LFInst_2_n2 ), .B(AddRoundKeyOutput[18]), .ZN(StateRegOutputF[14]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_4_LFInst_2_U3  ( .A(
        AddRoundKeyOutput[19]), .B(AddRoundKeyOutput[16]), .ZN(
        \StateRegOutputF_inst_LFInst_4_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_5_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst_LFInst_5_LFInst_0_n2 ), .B(AddRoundKeyOutput[21]), .ZN(StateRegOutputF[15]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_5_LFInst_0_U3  ( .A(
        AddRoundKeyOutput[22]), .B(AddRoundKeyOutput[20]), .ZN(
        \StateRegOutputF_inst_LFInst_5_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_5_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst_LFInst_5_LFInst_1_n2 ), .B(AddRoundKeyOutput[21]), .ZN(StateRegOutputF[16]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_5_LFInst_1_U3  ( .A(
        AddRoundKeyOutput[23]), .B(AddRoundKeyOutput[20]), .ZN(
        \StateRegOutputF_inst_LFInst_5_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_5_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst_LFInst_5_LFInst_2_n2 ), .B(AddRoundKeyOutput[22]), .ZN(StateRegOutputF[17]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_5_LFInst_2_U3  ( .A(
        AddRoundKeyOutput[23]), .B(AddRoundKeyOutput[20]), .ZN(
        \StateRegOutputF_inst_LFInst_5_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_6_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst_LFInst_6_LFInst_0_n2 ), .B(AddRoundKeyOutput[25]), .ZN(StateRegOutputF[18]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_6_LFInst_0_U3  ( .A(
        AddRoundKeyOutput[26]), .B(AddRoundKeyOutput[24]), .ZN(
        \StateRegOutputF_inst_LFInst_6_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_6_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst_LFInst_6_LFInst_1_n2 ), .B(AddRoundKeyOutput[25]), .ZN(StateRegOutputF[19]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_6_LFInst_1_U3  ( .A(
        AddRoundKeyOutput[27]), .B(AddRoundKeyOutput[24]), .ZN(
        \StateRegOutputF_inst_LFInst_6_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_6_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst_LFInst_6_LFInst_2_n2 ), .B(AddRoundKeyOutput[26]), .ZN(StateRegOutputF[20]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_6_LFInst_2_U3  ( .A(
        AddRoundKeyOutput[27]), .B(AddRoundKeyOutput[24]), .ZN(
        \StateRegOutputF_inst_LFInst_6_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_7_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst_LFInst_7_LFInst_0_n2 ), .B(AddRoundKeyOutput[29]), .ZN(StateRegOutputF[21]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_7_LFInst_0_U3  ( .A(
        AddRoundKeyOutput[30]), .B(AddRoundKeyOutput[28]), .ZN(
        \StateRegOutputF_inst_LFInst_7_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_7_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst_LFInst_7_LFInst_1_n2 ), .B(AddRoundKeyOutput[29]), .ZN(StateRegOutputF[22]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_7_LFInst_1_U3  ( .A(
        AddRoundKeyOutput[31]), .B(AddRoundKeyOutput[28]), .ZN(
        \StateRegOutputF_inst_LFInst_7_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_7_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst_LFInst_7_LFInst_2_n2 ), .B(AddRoundKeyOutput[30]), .ZN(StateRegOutputF[23]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_7_LFInst_2_U3  ( .A(
        AddRoundKeyOutput[31]), .B(AddRoundKeyOutput[28]), .ZN(
        \StateRegOutputF_inst_LFInst_7_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_8_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst_LFInst_8_LFInst_0_n2 ), .B(AddRoundKeyOutput[33]), .ZN(StateRegOutputF[24]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_8_LFInst_0_U3  ( .A(
        AddRoundKeyOutput[34]), .B(AddRoundKeyOutput[32]), .ZN(
        \StateRegOutputF_inst_LFInst_8_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_8_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst_LFInst_8_LFInst_1_n2 ), .B(AddRoundKeyOutput[33]), .ZN(StateRegOutputF[25]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_8_LFInst_1_U3  ( .A(
        AddRoundKeyOutput[35]), .B(AddRoundKeyOutput[32]), .ZN(
        \StateRegOutputF_inst_LFInst_8_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_8_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst_LFInst_8_LFInst_2_n2 ), .B(AddRoundKeyOutput[34]), .ZN(StateRegOutputF[26]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_8_LFInst_2_U3  ( .A(
        AddRoundKeyOutput[35]), .B(AddRoundKeyOutput[32]), .ZN(
        \StateRegOutputF_inst_LFInst_8_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_9_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst_LFInst_9_LFInst_0_n2 ), .B(AddRoundKeyOutput[37]), .ZN(StateRegOutputF[27]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_9_LFInst_0_U3  ( .A(
        AddRoundKeyOutput[38]), .B(AddRoundKeyOutput[36]), .ZN(
        \StateRegOutputF_inst_LFInst_9_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_9_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst_LFInst_9_LFInst_1_n2 ), .B(AddRoundKeyOutput[37]), .ZN(StateRegOutputF[28]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_9_LFInst_1_U3  ( .A(
        AddRoundKeyOutput[39]), .B(AddRoundKeyOutput[36]), .ZN(
        \StateRegOutputF_inst_LFInst_9_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_9_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst_LFInst_9_LFInst_2_n2 ), .B(AddRoundKeyOutput[38]), .ZN(StateRegOutputF[29]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_9_LFInst_2_U3  ( .A(
        AddRoundKeyOutput[39]), .B(AddRoundKeyOutput[36]), .ZN(
        \StateRegOutputF_inst_LFInst_9_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_10_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst_LFInst_10_LFInst_0_n2 ), .B(
        AddRoundKeyOutput[41]), .ZN(StateRegOutputF[30]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_10_LFInst_0_U3  ( .A(
        AddRoundKeyOutput[42]), .B(AddRoundKeyOutput[40]), .ZN(
        \StateRegOutputF_inst_LFInst_10_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_10_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst_LFInst_10_LFInst_1_n2 ), .B(
        AddRoundKeyOutput[41]), .ZN(StateRegOutputF[31]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_10_LFInst_1_U3  ( .A(
        AddRoundKeyOutput[43]), .B(AddRoundKeyOutput[40]), .ZN(
        \StateRegOutputF_inst_LFInst_10_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_10_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst_LFInst_10_LFInst_2_n2 ), .B(
        AddRoundKeyOutput[42]), .ZN(StateRegOutputF[32]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_10_LFInst_2_U3  ( .A(
        AddRoundKeyOutput[43]), .B(AddRoundKeyOutput[40]), .ZN(
        \StateRegOutputF_inst_LFInst_10_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_11_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst_LFInst_11_LFInst_0_n2 ), .B(
        AddRoundKeyOutput[45]), .ZN(StateRegOutputF[33]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_11_LFInst_0_U3  ( .A(
        AddRoundKeyOutput[46]), .B(AddRoundKeyOutput[44]), .ZN(
        \StateRegOutputF_inst_LFInst_11_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_11_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst_LFInst_11_LFInst_1_n2 ), .B(
        AddRoundKeyOutput[45]), .ZN(StateRegOutputF[34]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_11_LFInst_1_U3  ( .A(
        AddRoundKeyOutput[47]), .B(AddRoundKeyOutput[44]), .ZN(
        \StateRegOutputF_inst_LFInst_11_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_11_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst_LFInst_11_LFInst_2_n2 ), .B(
        AddRoundKeyOutput[46]), .ZN(StateRegOutputF[35]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_11_LFInst_2_U3  ( .A(
        AddRoundKeyOutput[47]), .B(AddRoundKeyOutput[44]), .ZN(
        \StateRegOutputF_inst_LFInst_11_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_12_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst_LFInst_12_LFInst_0_n2 ), .B(
        AddRoundKeyOutput[49]), .ZN(StateRegOutputF[36]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_12_LFInst_0_U3  ( .A(
        AddRoundKeyOutput[50]), .B(AddRoundKeyOutput[48]), .ZN(
        \StateRegOutputF_inst_LFInst_12_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_12_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst_LFInst_12_LFInst_1_n2 ), .B(
        AddRoundKeyOutput[49]), .ZN(StateRegOutputF[37]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_12_LFInst_1_U3  ( .A(
        AddRoundKeyOutput[51]), .B(AddRoundKeyOutput[48]), .ZN(
        \StateRegOutputF_inst_LFInst_12_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_12_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst_LFInst_12_LFInst_2_n2 ), .B(
        AddRoundKeyOutput[50]), .ZN(StateRegOutputF[38]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_12_LFInst_2_U3  ( .A(
        AddRoundKeyOutput[51]), .B(AddRoundKeyOutput[48]), .ZN(
        \StateRegOutputF_inst_LFInst_12_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_13_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst_LFInst_13_LFInst_0_n2 ), .B(
        AddRoundKeyOutput[53]), .ZN(StateRegOutputF[39]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_13_LFInst_0_U3  ( .A(
        AddRoundKeyOutput[54]), .B(AddRoundKeyOutput[52]), .ZN(
        \StateRegOutputF_inst_LFInst_13_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_13_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst_LFInst_13_LFInst_1_n2 ), .B(
        AddRoundKeyOutput[53]), .ZN(StateRegOutputF[40]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_13_LFInst_1_U3  ( .A(
        AddRoundKeyOutput[55]), .B(AddRoundKeyOutput[52]), .ZN(
        \StateRegOutputF_inst_LFInst_13_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_13_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst_LFInst_13_LFInst_2_n2 ), .B(
        AddRoundKeyOutput[54]), .ZN(StateRegOutputF[41]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_13_LFInst_2_U3  ( .A(
        AddRoundKeyOutput[55]), .B(AddRoundKeyOutput[52]), .ZN(
        \StateRegOutputF_inst_LFInst_13_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_14_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst_LFInst_14_LFInst_0_n2 ), .B(
        AddRoundKeyOutput[57]), .ZN(StateRegOutputF[42]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_14_LFInst_0_U3  ( .A(
        AddRoundKeyOutput[58]), .B(AddRoundKeyOutput[56]), .ZN(
        \StateRegOutputF_inst_LFInst_14_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_14_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst_LFInst_14_LFInst_1_n2 ), .B(
        AddRoundKeyOutput[57]), .ZN(StateRegOutputF[43]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_14_LFInst_1_U3  ( .A(
        AddRoundKeyOutput[59]), .B(AddRoundKeyOutput[56]), .ZN(
        \StateRegOutputF_inst_LFInst_14_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_14_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst_LFInst_14_LFInst_2_n2 ), .B(
        AddRoundKeyOutput[58]), .ZN(StateRegOutputF[44]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_14_LFInst_2_U3  ( .A(
        AddRoundKeyOutput[59]), .B(AddRoundKeyOutput[56]), .ZN(
        \StateRegOutputF_inst_LFInst_14_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_15_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst_LFInst_15_LFInst_0_n2 ), .B(
        AddRoundKeyOutput[61]), .ZN(StateRegOutputF[45]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_15_LFInst_0_U3  ( .A(
        AddRoundKeyOutput[62]), .B(AddRoundKeyOutput[60]), .ZN(
        \StateRegOutputF_inst_LFInst_15_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_15_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst_LFInst_15_LFInst_1_n2 ), .B(
        AddRoundKeyOutput[61]), .ZN(StateRegOutputF[46]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_15_LFInst_1_U3  ( .A(
        AddRoundKeyOutput[63]), .B(AddRoundKeyOutput[60]), .ZN(
        \StateRegOutputF_inst_LFInst_15_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_15_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst_LFInst_15_LFInst_2_n2 ), .B(
        AddRoundKeyOutput[62]), .ZN(StateRegOutputF[47]) );
  XNOR2_X1 \StateRegOutputF_inst_LFInst_15_LFInst_2_U3  ( .A(
        AddRoundKeyOutput[63]), .B(AddRoundKeyOutput[60]), .ZN(
        \StateRegOutputF_inst_LFInst_15_LFInst_2_n2 ) );
  INV_X1 \CipherErrorVecGen_XORInst_0_0_U2  ( .A(
        \CipherErrorVecGen_XORInst_0_0_n4 ), .ZN(CipherErrorVec[0]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_0_0_U1  ( .A(StateRegOutputF[0]), .B(
        Red_AddRoundKeyOutput[0]), .ZN(\CipherErrorVecGen_XORInst_0_0_n4 ) );
  INV_X1 \CipherErrorVecGen_XORInst_0_1_U2  ( .A(
        \CipherErrorVecGen_XORInst_0_1_n2 ), .ZN(CipherErrorVec[1]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_0_1_U1  ( .A(StateRegOutputF[1]), .B(
        Red_AddRoundKeyOutput[1]), .ZN(\CipherErrorVecGen_XORInst_0_1_n2 ) );
  INV_X1 \CipherErrorVecGen_XORInst_0_2_U2  ( .A(
        \CipherErrorVecGen_XORInst_0_2_n3 ), .ZN(CipherErrorVec[2]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_0_2_U1  ( .A(StateRegOutputF[2]), .B(
        Red_AddRoundKeyOutput[2]), .ZN(\CipherErrorVecGen_XORInst_0_2_n3 ) );
  INV_X1 \CipherErrorVecGen_XORInst_1_0_U2  ( .A(
        \CipherErrorVecGen_XORInst_1_0_n4 ), .ZN(CipherErrorVec[3]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_1_0_U1  ( .A(StateRegOutputF[3]), .B(
        Red_AddRoundKeyOutput[3]), .ZN(\CipherErrorVecGen_XORInst_1_0_n4 ) );
  INV_X1 \CipherErrorVecGen_XORInst_1_1_U2  ( .A(
        \CipherErrorVecGen_XORInst_1_1_n2 ), .ZN(CipherErrorVec[4]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_1_1_U1  ( .A(StateRegOutputF[4]), .B(
        Red_AddRoundKeyOutput[4]), .ZN(\CipherErrorVecGen_XORInst_1_1_n2 ) );
  INV_X1 \CipherErrorVecGen_XORInst_1_2_U2  ( .A(
        \CipherErrorVecGen_XORInst_1_2_n3 ), .ZN(CipherErrorVec[5]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_1_2_U1  ( .A(StateRegOutputF[5]), .B(
        Red_AddRoundKeyOutput[5]), .ZN(\CipherErrorVecGen_XORInst_1_2_n3 ) );
  INV_X1 \CipherErrorVecGen_XORInst_2_0_U2  ( .A(
        \CipherErrorVecGen_XORInst_2_0_n4 ), .ZN(CipherErrorVec[6]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_2_0_U1  ( .A(StateRegOutputF[6]), .B(
        Red_AddRoundKeyOutput[6]), .ZN(\CipherErrorVecGen_XORInst_2_0_n4 ) );
  INV_X1 \CipherErrorVecGen_XORInst_2_1_U2  ( .A(
        \CipherErrorVecGen_XORInst_2_1_n2 ), .ZN(CipherErrorVec[7]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_2_1_U1  ( .A(StateRegOutputF[7]), .B(
        Red_AddRoundKeyOutput[7]), .ZN(\CipherErrorVecGen_XORInst_2_1_n2 ) );
  INV_X1 \CipherErrorVecGen_XORInst_2_2_U2  ( .A(
        \CipherErrorVecGen_XORInst_2_2_n3 ), .ZN(CipherErrorVec[8]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_2_2_U1  ( .A(StateRegOutputF[8]), .B(
        Red_AddRoundKeyOutput[8]), .ZN(\CipherErrorVecGen_XORInst_2_2_n3 ) );
  INV_X1 \CipherErrorVecGen_XORInst_3_0_U2  ( .A(
        \CipherErrorVecGen_XORInst_3_0_n4 ), .ZN(CipherErrorVec[9]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_3_0_U1  ( .A(StateRegOutputF[9]), .B(
        Red_AddRoundKeyOutput[9]), .ZN(\CipherErrorVecGen_XORInst_3_0_n4 ) );
  INV_X1 \CipherErrorVecGen_XORInst_3_1_U2  ( .A(
        \CipherErrorVecGen_XORInst_3_1_n2 ), .ZN(CipherErrorVec[10]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_3_1_U1  ( .A(StateRegOutputF[10]), .B(
        Red_AddRoundKeyOutput[10]), .ZN(\CipherErrorVecGen_XORInst_3_1_n2 ) );
  INV_X1 \CipherErrorVecGen_XORInst_3_2_U2  ( .A(
        \CipherErrorVecGen_XORInst_3_2_n3 ), .ZN(CipherErrorVec[11]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_3_2_U1  ( .A(StateRegOutputF[11]), .B(
        Red_AddRoundKeyOutput[11]), .ZN(\CipherErrorVecGen_XORInst_3_2_n3 ) );
  INV_X1 \CipherErrorVecGen_XORInst_4_0_U2  ( .A(
        \CipherErrorVecGen_XORInst_4_0_n4 ), .ZN(CipherErrorVec[12]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_4_0_U1  ( .A(StateRegOutputF[12]), .B(
        Red_AddRoundKeyOutput[12]), .ZN(\CipherErrorVecGen_XORInst_4_0_n4 ) );
  INV_X1 \CipherErrorVecGen_XORInst_4_1_U2  ( .A(
        \CipherErrorVecGen_XORInst_4_1_n2 ), .ZN(CipherErrorVec[13]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_4_1_U1  ( .A(StateRegOutputF[13]), .B(
        Red_AddRoundKeyOutput[13]), .ZN(\CipherErrorVecGen_XORInst_4_1_n2 ) );
  INV_X1 \CipherErrorVecGen_XORInst_4_2_U2  ( .A(
        \CipherErrorVecGen_XORInst_4_2_n3 ), .ZN(CipherErrorVec[14]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_4_2_U1  ( .A(StateRegOutputF[14]), .B(
        Red_AddRoundKeyOutput[14]), .ZN(\CipherErrorVecGen_XORInst_4_2_n3 ) );
  INV_X1 \CipherErrorVecGen_XORInst_5_0_U2  ( .A(
        \CipherErrorVecGen_XORInst_5_0_n4 ), .ZN(CipherErrorVec[15]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_5_0_U1  ( .A(StateRegOutputF[15]), .B(
        Red_AddRoundKeyOutput[15]), .ZN(\CipherErrorVecGen_XORInst_5_0_n4 ) );
  INV_X1 \CipherErrorVecGen_XORInst_5_1_U2  ( .A(
        \CipherErrorVecGen_XORInst_5_1_n2 ), .ZN(CipherErrorVec[16]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_5_1_U1  ( .A(StateRegOutputF[16]), .B(
        Red_AddRoundKeyOutput[16]), .ZN(\CipherErrorVecGen_XORInst_5_1_n2 ) );
  INV_X1 \CipherErrorVecGen_XORInst_5_2_U2  ( .A(
        \CipherErrorVecGen_XORInst_5_2_n3 ), .ZN(CipherErrorVec[17]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_5_2_U1  ( .A(StateRegOutputF[17]), .B(
        Red_AddRoundKeyOutput[17]), .ZN(\CipherErrorVecGen_XORInst_5_2_n3 ) );
  INV_X1 \CipherErrorVecGen_XORInst_6_0_U2  ( .A(
        \CipherErrorVecGen_XORInst_6_0_n4 ), .ZN(CipherErrorVec[18]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_6_0_U1  ( .A(StateRegOutputF[18]), .B(
        Red_AddRoundKeyOutput[18]), .ZN(\CipherErrorVecGen_XORInst_6_0_n4 ) );
  INV_X1 \CipherErrorVecGen_XORInst_6_1_U2  ( .A(
        \CipherErrorVecGen_XORInst_6_1_n2 ), .ZN(CipherErrorVec[19]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_6_1_U1  ( .A(StateRegOutputF[19]), .B(
        Red_AddRoundKeyOutput[19]), .ZN(\CipherErrorVecGen_XORInst_6_1_n2 ) );
  INV_X1 \CipherErrorVecGen_XORInst_6_2_U2  ( .A(
        \CipherErrorVecGen_XORInst_6_2_n3 ), .ZN(CipherErrorVec[20]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_6_2_U1  ( .A(StateRegOutputF[20]), .B(
        Red_AddRoundKeyOutput[20]), .ZN(\CipherErrorVecGen_XORInst_6_2_n3 ) );
  INV_X1 \CipherErrorVecGen_XORInst_7_0_U2  ( .A(
        \CipherErrorVecGen_XORInst_7_0_n4 ), .ZN(CipherErrorVec[21]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_7_0_U1  ( .A(StateRegOutputF[21]), .B(
        Red_AddRoundKeyOutput[21]), .ZN(\CipherErrorVecGen_XORInst_7_0_n4 ) );
  INV_X1 \CipherErrorVecGen_XORInst_7_1_U2  ( .A(
        \CipherErrorVecGen_XORInst_7_1_n2 ), .ZN(CipherErrorVec[22]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_7_1_U1  ( .A(StateRegOutputF[22]), .B(
        Red_AddRoundKeyOutput[22]), .ZN(\CipherErrorVecGen_XORInst_7_1_n2 ) );
  INV_X1 \CipherErrorVecGen_XORInst_7_2_U2  ( .A(
        \CipherErrorVecGen_XORInst_7_2_n3 ), .ZN(CipherErrorVec[23]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_7_2_U1  ( .A(StateRegOutputF[23]), .B(
        Red_AddRoundKeyOutput[23]), .ZN(\CipherErrorVecGen_XORInst_7_2_n3 ) );
  INV_X1 \CipherErrorVecGen_XORInst_8_0_U2  ( .A(
        \CipherErrorVecGen_XORInst_8_0_n4 ), .ZN(CipherErrorVec[24]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_8_0_U1  ( .A(StateRegOutputF[24]), .B(
        Red_AddRoundKeyOutput[24]), .ZN(\CipherErrorVecGen_XORInst_8_0_n4 ) );
  INV_X1 \CipherErrorVecGen_XORInst_8_1_U2  ( .A(
        \CipherErrorVecGen_XORInst_8_1_n2 ), .ZN(CipherErrorVec[25]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_8_1_U1  ( .A(StateRegOutputF[25]), .B(
        Red_AddRoundKeyOutput[25]), .ZN(\CipherErrorVecGen_XORInst_8_1_n2 ) );
  INV_X1 \CipherErrorVecGen_XORInst_8_2_U2  ( .A(
        \CipherErrorVecGen_XORInst_8_2_n3 ), .ZN(CipherErrorVec[26]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_8_2_U1  ( .A(StateRegOutputF[26]), .B(
        Red_AddRoundKeyOutput[26]), .ZN(\CipherErrorVecGen_XORInst_8_2_n3 ) );
  INV_X1 \CipherErrorVecGen_XORInst_9_0_U2  ( .A(
        \CipherErrorVecGen_XORInst_9_0_n4 ), .ZN(CipherErrorVec[27]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_9_0_U1  ( .A(StateRegOutputF[27]), .B(
        Red_AddRoundKeyOutput[27]), .ZN(\CipherErrorVecGen_XORInst_9_0_n4 ) );
  INV_X1 \CipherErrorVecGen_XORInst_9_1_U2  ( .A(
        \CipherErrorVecGen_XORInst_9_1_n2 ), .ZN(CipherErrorVec[28]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_9_1_U1  ( .A(StateRegOutputF[28]), .B(
        Red_AddRoundKeyOutput[28]), .ZN(\CipherErrorVecGen_XORInst_9_1_n2 ) );
  INV_X1 \CipherErrorVecGen_XORInst_9_2_U2  ( .A(
        \CipherErrorVecGen_XORInst_9_2_n3 ), .ZN(CipherErrorVec[29]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_9_2_U1  ( .A(StateRegOutputF[29]), .B(
        Red_AddRoundKeyOutput[29]), .ZN(\CipherErrorVecGen_XORInst_9_2_n3 ) );
  INV_X1 \CipherErrorVecGen_XORInst_10_0_U2  ( .A(
        \CipherErrorVecGen_XORInst_10_0_n4 ), .ZN(CipherErrorVec[30]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_10_0_U1  ( .A(StateRegOutputF[30]), .B(
        Red_AddRoundKeyOutput[30]), .ZN(\CipherErrorVecGen_XORInst_10_0_n4 )
         );
  INV_X1 \CipherErrorVecGen_XORInst_10_1_U2  ( .A(
        \CipherErrorVecGen_XORInst_10_1_n2 ), .ZN(CipherErrorVec[31]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_10_1_U1  ( .A(StateRegOutputF[31]), .B(
        Red_AddRoundKeyOutput[31]), .ZN(\CipherErrorVecGen_XORInst_10_1_n2 )
         );
  INV_X1 \CipherErrorVecGen_XORInst_10_2_U2  ( .A(
        \CipherErrorVecGen_XORInst_10_2_n3 ), .ZN(CipherErrorVec[32]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_10_2_U1  ( .A(StateRegOutputF[32]), .B(
        Red_AddRoundKeyOutput[32]), .ZN(\CipherErrorVecGen_XORInst_10_2_n3 )
         );
  INV_X1 \CipherErrorVecGen_XORInst_11_0_U2  ( .A(
        \CipherErrorVecGen_XORInst_11_0_n4 ), .ZN(CipherErrorVec[33]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_11_0_U1  ( .A(StateRegOutputF[33]), .B(
        Red_AddRoundKeyOutput[33]), .ZN(\CipherErrorVecGen_XORInst_11_0_n4 )
         );
  INV_X1 \CipherErrorVecGen_XORInst_11_1_U2  ( .A(
        \CipherErrorVecGen_XORInst_11_1_n2 ), .ZN(CipherErrorVec[34]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_11_1_U1  ( .A(StateRegOutputF[34]), .B(
        Red_AddRoundKeyOutput[34]), .ZN(\CipherErrorVecGen_XORInst_11_1_n2 )
         );
  INV_X1 \CipherErrorVecGen_XORInst_11_2_U2  ( .A(
        \CipherErrorVecGen_XORInst_11_2_n3 ), .ZN(CipherErrorVec[35]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_11_2_U1  ( .A(StateRegOutputF[35]), .B(
        Red_AddRoundKeyOutput[35]), .ZN(\CipherErrorVecGen_XORInst_11_2_n3 )
         );
  INV_X1 \CipherErrorVecGen_XORInst_12_0_U2  ( .A(
        \CipherErrorVecGen_XORInst_12_0_n4 ), .ZN(CipherErrorVec[36]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_12_0_U1  ( .A(StateRegOutputF[36]), .B(
        Red_AddRoundKeyOutput[36]), .ZN(\CipherErrorVecGen_XORInst_12_0_n4 )
         );
  INV_X1 \CipherErrorVecGen_XORInst_12_1_U2  ( .A(
        \CipherErrorVecGen_XORInst_12_1_n2 ), .ZN(CipherErrorVec[37]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_12_1_U1  ( .A(StateRegOutputF[37]), .B(
        Red_AddRoundKeyOutput[37]), .ZN(\CipherErrorVecGen_XORInst_12_1_n2 )
         );
  INV_X1 \CipherErrorVecGen_XORInst_12_2_U2  ( .A(
        \CipherErrorVecGen_XORInst_12_2_n3 ), .ZN(CipherErrorVec[38]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_12_2_U1  ( .A(StateRegOutputF[38]), .B(
        Red_AddRoundKeyOutput[38]), .ZN(\CipherErrorVecGen_XORInst_12_2_n3 )
         );
  INV_X1 \CipherErrorVecGen_XORInst_13_0_U2  ( .A(
        \CipherErrorVecGen_XORInst_13_0_n4 ), .ZN(CipherErrorVec[39]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_13_0_U1  ( .A(StateRegOutputF[39]), .B(
        Red_AddRoundKeyOutput[39]), .ZN(\CipherErrorVecGen_XORInst_13_0_n4 )
         );
  INV_X1 \CipherErrorVecGen_XORInst_13_1_U2  ( .A(
        \CipherErrorVecGen_XORInst_13_1_n2 ), .ZN(CipherErrorVec[40]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_13_1_U1  ( .A(StateRegOutputF[40]), .B(
        Red_AddRoundKeyOutput[40]), .ZN(\CipherErrorVecGen_XORInst_13_1_n2 )
         );
  INV_X1 \CipherErrorVecGen_XORInst_13_2_U2  ( .A(
        \CipherErrorVecGen_XORInst_13_2_n3 ), .ZN(CipherErrorVec[41]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_13_2_U1  ( .A(StateRegOutputF[41]), .B(
        Red_AddRoundKeyOutput[41]), .ZN(\CipherErrorVecGen_XORInst_13_2_n3 )
         );
  INV_X1 \CipherErrorVecGen_XORInst_14_0_U2  ( .A(
        \CipherErrorVecGen_XORInst_14_0_n4 ), .ZN(CipherErrorVec[42]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_14_0_U1  ( .A(StateRegOutputF[42]), .B(
        Red_AddRoundKeyOutput[42]), .ZN(\CipherErrorVecGen_XORInst_14_0_n4 )
         );
  INV_X1 \CipherErrorVecGen_XORInst_14_1_U2  ( .A(
        \CipherErrorVecGen_XORInst_14_1_n2 ), .ZN(CipherErrorVec[43]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_14_1_U1  ( .A(StateRegOutputF[43]), .B(
        Red_AddRoundKeyOutput[43]), .ZN(\CipherErrorVecGen_XORInst_14_1_n2 )
         );
  INV_X1 \CipherErrorVecGen_XORInst_14_2_U2  ( .A(
        \CipherErrorVecGen_XORInst_14_2_n3 ), .ZN(CipherErrorVec[44]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_14_2_U1  ( .A(StateRegOutputF[44]), .B(
        Red_AddRoundKeyOutput[44]), .ZN(\CipherErrorVecGen_XORInst_14_2_n3 )
         );
  INV_X1 \CipherErrorVecGen_XORInst_15_0_U2  ( .A(
        \CipherErrorVecGen_XORInst_15_0_n4 ), .ZN(CipherErrorVec[45]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_15_0_U1  ( .A(StateRegOutputF[45]), .B(
        Red_AddRoundKeyOutput[45]), .ZN(\CipherErrorVecGen_XORInst_15_0_n4 )
         );
  INV_X1 \CipherErrorVecGen_XORInst_15_1_U2  ( .A(
        \CipherErrorVecGen_XORInst_15_1_n2 ), .ZN(CipherErrorVec[46]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_15_1_U1  ( .A(StateRegOutputF[46]), .B(
        Red_AddRoundKeyOutput[46]), .ZN(\CipherErrorVecGen_XORInst_15_1_n2 )
         );
  INV_X1 \CipherErrorVecGen_XORInst_15_2_U2  ( .A(
        \CipherErrorVecGen_XORInst_15_2_n3 ), .ZN(CipherErrorVec[47]) );
  XNOR2_X1 \CipherErrorVecGen_XORInst_15_2_U1  ( .A(StateRegOutputF[47]), .B(
        Red_AddRoundKeyOutput[47]), .ZN(\CipherErrorVecGen_XORInst_15_2_n3 )
         );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n35 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n34 ), .ZN(
        Red_PermutationInput[0]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U18  ( .A1(
        CipherErrorVec[2]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n33 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n34 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U17  ( .A1(
        CipherErrorVec[0]), .A2(CipherErrorVec[1]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n32 ), .B(
        AddRoundKeyOutput[1]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n30 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U13  ( .A(
        AddRoundKeyOutput[0]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n28 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U12  ( .A1(
        CipherErrorVec[1]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n26 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n27 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U11  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U10  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n24 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n23 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n31 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n23 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U8  ( .A(
        AddRoundKeyOutput[3]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n22 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U7  ( .A1(
        CipherErrorVec[0]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n21 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n22 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U6  ( .A1(
        CipherErrorVec[1]), .A2(CipherErrorVec[2]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U5  ( .A(
        AddRoundKeyOutput[2]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n20 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U4  ( .A1(
        CipherErrorVec[1]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n25 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U3  ( .A1(
        CipherErrorVec[2]), .A2(CipherErrorVec[0]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n25 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U22  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n36 ), .ZN(
        Red_PermutationInput[1]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n36 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n33 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n34 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U18  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n30 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n37 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U17  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n29 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n28 ), .B(
        AddRoundKeyOutput[0]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n31 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n28 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U14  ( .A(
        AddRoundKeyOutput[2]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n25 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n35 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U13  ( .A1(
        CipherErrorVec[1]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n24 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U12  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n23 ), .A2(CipherErrorVec[2]), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n32 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n22 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n30 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U10  ( .A(
        AddRoundKeyOutput[3]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n21 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n22 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U9  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n23 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n21 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U8  ( .A1(
        CipherErrorVec[1]), .A2(CipherErrorVec[2]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n27 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U7  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n20 ), .B(
        AddRoundKeyOutput[1]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n32 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U6  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n19 ), .A2(CipherErrorVec[2]), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U5  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n23 ), .A2(CipherErrorVec[1]), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n19 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U4  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U3  ( .A(CipherErrorVec[0]), 
        .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n36 ), .ZN(
        Red_PermutationInput[2]) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n36 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U19  ( .A(
        AddRoundKeyOutput[1]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n33 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n34 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U18  ( .A1(
        CipherErrorVec[2]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n32 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n33 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U17  ( .A1(
        CipherErrorVec[0]), .A2(CipherErrorVec[1]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U16  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n31 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n37 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U13  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n26 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U12  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n25 ), .B(
        AddRoundKeyOutput[2]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n28 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n24 ), .A2(CipherErrorVec[1]), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U10  ( .A1(
        CipherErrorVec[0]), .A2(CipherErrorVec[2]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n24 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n29 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n30 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n27 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U8  ( .A(
        AddRoundKeyOutput[0]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n23 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n30 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U7  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n22 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U6  ( .A(CipherErrorVec[0]), 
        .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n22 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U5  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n20 ), .B(
        AddRoundKeyOutput[3]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U4  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n21 ), .A2(CipherErrorVec[0]), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U3  ( .A1(
        CipherErrorVec[1]), .A2(CipherErrorVec[2]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n35 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n34 ), .ZN(
        Red_PermutationInput[3]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U18  ( .A1(
        CipherErrorVec[5]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n33 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n34 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U17  ( .A1(
        CipherErrorVec[3]), .A2(CipherErrorVec[4]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n32 ), .B(
        AddRoundKeyOutput[5]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n30 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U13  ( .A(
        AddRoundKeyOutput[4]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n28 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U12  ( .A1(
        CipherErrorVec[4]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n26 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n27 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U11  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U10  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n24 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n23 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n31 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n23 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U8  ( .A(
        AddRoundKeyOutput[7]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n22 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U7  ( .A1(
        CipherErrorVec[3]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n21 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n22 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U6  ( .A1(
        CipherErrorVec[4]), .A2(CipherErrorVec[5]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U5  ( .A(
        AddRoundKeyOutput[6]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n20 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U4  ( .A1(
        CipherErrorVec[4]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n25 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U3  ( .A1(
        CipherErrorVec[5]), .A2(CipherErrorVec[3]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n25 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U22  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n36 ), .ZN(
        Red_PermutationInput[4]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n36 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n33 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n34 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U18  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n30 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n37 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U17  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n29 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n28 ), .B(
        AddRoundKeyOutput[4]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n31 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n28 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U14  ( .A(
        AddRoundKeyOutput[6]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n25 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n35 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U13  ( .A1(
        CipherErrorVec[4]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n24 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U12  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n23 ), .A2(CipherErrorVec[5]), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n32 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n22 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n30 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U10  ( .A(
        AddRoundKeyOutput[7]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n21 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n22 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U9  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n23 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n21 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U8  ( .A1(
        CipherErrorVec[4]), .A2(CipherErrorVec[5]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n27 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U7  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n20 ), .B(
        AddRoundKeyOutput[5]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n32 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U6  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n19 ), .A2(CipherErrorVec[5]), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U5  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n23 ), .A2(CipherErrorVec[4]), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n19 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U4  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U3  ( .A(CipherErrorVec[3]), 
        .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n36 ), .ZN(
        Red_PermutationInput[5]) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n36 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U19  ( .A(
        AddRoundKeyOutput[5]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n33 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n34 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U18  ( .A1(
        CipherErrorVec[5]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n32 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n33 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U17  ( .A1(
        CipherErrorVec[3]), .A2(CipherErrorVec[4]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U16  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n31 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n37 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U13  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n26 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U12  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n25 ), .B(
        AddRoundKeyOutput[6]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n28 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n24 ), .A2(CipherErrorVec[4]), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U10  ( .A1(
        CipherErrorVec[3]), .A2(CipherErrorVec[5]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n24 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n29 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n30 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n27 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U8  ( .A(
        AddRoundKeyOutput[4]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n23 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n30 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U7  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n22 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U6  ( .A(CipherErrorVec[3]), 
        .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n22 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U5  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n20 ), .B(
        AddRoundKeyOutput[7]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U4  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n21 ), .A2(CipherErrorVec[3]), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U3  ( .A1(
        CipherErrorVec[4]), .A2(CipherErrorVec[5]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n35 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n34 ), .ZN(
        Red_PermutationInput[6]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U18  ( .A1(
        CipherErrorVec[8]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n33 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n34 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U17  ( .A1(
        CipherErrorVec[6]), .A2(CipherErrorVec[7]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n32 ), .B(
        AddRoundKeyOutput[9]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n30 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U13  ( .A(
        AddRoundKeyOutput[8]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n28 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U12  ( .A1(
        CipherErrorVec[7]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n26 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n27 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U11  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U10  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n24 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n23 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n31 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n23 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U8  ( .A(
        AddRoundKeyOutput[11]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n22 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U7  ( .A1(
        CipherErrorVec[6]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n21 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n22 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U6  ( .A1(
        CipherErrorVec[7]), .A2(CipherErrorVec[8]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U5  ( .A(
        AddRoundKeyOutput[10]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n20 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U4  ( .A1(
        CipherErrorVec[7]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n25 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U3  ( .A1(
        CipherErrorVec[8]), .A2(CipherErrorVec[6]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n25 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U22  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n36 ), .ZN(
        Red_PermutationInput[7]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n36 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n33 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n34 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U18  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n30 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n37 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U17  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n29 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n28 ), .B(
        AddRoundKeyOutput[8]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n31 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n28 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U14  ( .A(
        AddRoundKeyOutput[10]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n25 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n35 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U13  ( .A1(
        CipherErrorVec[7]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n24 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U12  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n23 ), .A2(CipherErrorVec[8]), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n32 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n22 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n30 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U10  ( .A(
        AddRoundKeyOutput[11]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n21 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n22 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U9  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n23 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n21 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U8  ( .A1(
        CipherErrorVec[7]), .A2(CipherErrorVec[8]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n27 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U7  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n20 ), .B(
        AddRoundKeyOutput[9]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n32 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U6  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n19 ), .A2(CipherErrorVec[8]), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U5  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n23 ), .A2(CipherErrorVec[7]), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n19 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U4  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U3  ( .A(CipherErrorVec[6]), 
        .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n36 ), .ZN(
        Red_PermutationInput[8]) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n36 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U19  ( .A(
        AddRoundKeyOutput[9]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n33 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n34 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U18  ( .A1(
        CipherErrorVec[8]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n32 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n33 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U17  ( .A1(
        CipherErrorVec[6]), .A2(CipherErrorVec[7]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U16  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n31 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n37 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U13  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n26 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U12  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n25 ), .B(
        AddRoundKeyOutput[10]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n28 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n24 ), .A2(CipherErrorVec[7]), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U10  ( .A1(
        CipherErrorVec[6]), .A2(CipherErrorVec[8]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n24 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n29 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n30 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n27 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U8  ( .A(
        AddRoundKeyOutput[8]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n23 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n30 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U7  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n22 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U6  ( .A(CipherErrorVec[6]), 
        .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n22 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U5  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n20 ), .B(
        AddRoundKeyOutput[11]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U4  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n21 ), .A2(CipherErrorVec[6]), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U3  ( .A1(
        CipherErrorVec[7]), .A2(CipherErrorVec[8]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n35 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n34 ), .ZN(
        Red_PermutationInput[9]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U18  ( .A1(
        CipherErrorVec[11]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n33 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n34 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U17  ( .A1(
        CipherErrorVec[9]), .A2(CipherErrorVec[10]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n32 ), .B(
        AddRoundKeyOutput[13]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n30 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U13  ( .A(
        AddRoundKeyOutput[12]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n28 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U12  ( .A1(
        CipherErrorVec[10]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n27 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U11  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U10  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n24 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n23 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n31 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n23 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U8  ( .A(
        AddRoundKeyOutput[15]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n22 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U7  ( .A1(
        CipherErrorVec[9]), .A2(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n21 ), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n22 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U6  ( .A1(
        CipherErrorVec[10]), .A2(CipherErrorVec[11]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U5  ( .A(
        AddRoundKeyOutput[14]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n20 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U4  ( .A1(
        CipherErrorVec[10]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U3  ( .A1(
        CipherErrorVec[11]), .A2(CipherErrorVec[9]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n25 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U22  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n36 ), .ZN(
        Red_PermutationInput[10]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n36 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n33 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n34 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U18  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n30 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n37 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U17  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n29 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n28 ), .B(
        AddRoundKeyOutput[12]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n31 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n28 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U14  ( .A(
        AddRoundKeyOutput[14]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n25 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n35 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U13  ( .A1(
        CipherErrorVec[10]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n24 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U12  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n23 ), .A2(
        CipherErrorVec[11]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n32 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n22 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n30 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U10  ( .A(
        AddRoundKeyOutput[15]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n21 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n22 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U9  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n23 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n21 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U8  ( .A1(
        CipherErrorVec[10]), .A2(CipherErrorVec[11]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n27 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U7  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n20 ), .B(
        AddRoundKeyOutput[13]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n32 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U6  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n19 ), .A2(
        CipherErrorVec[11]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U5  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n23 ), .A2(
        CipherErrorVec[10]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n19 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U4  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U3  ( .A(CipherErrorVec[9]), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n36 ), .ZN(
        Red_PermutationInput[11]) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n36 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U19  ( .A(
        AddRoundKeyOutput[13]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n33 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n34 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U18  ( .A1(
        CipherErrorVec[11]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n33 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U17  ( .A1(
        CipherErrorVec[9]), .A2(CipherErrorVec[10]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U16  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n31 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n37 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U13  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n26 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U12  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n25 ), .B(
        AddRoundKeyOutput[14]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n28 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n24 ), .A2(
        CipherErrorVec[10]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U10  ( .A1(
        CipherErrorVec[9]), .A2(CipherErrorVec[11]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n24 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n29 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n30 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n27 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U8  ( .A(
        AddRoundKeyOutput[12]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n23 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n30 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U7  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n22 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U6  ( .A(CipherErrorVec[9]), .ZN(\SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n22 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U5  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n20 ), .B(
        AddRoundKeyOutput[15]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U4  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n21 ), .A2(
        CipherErrorVec[9]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U3  ( .A1(
        CipherErrorVec[10]), .A2(CipherErrorVec[11]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n35 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n34 ), .ZN(
        Red_PermutationInput[12]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U18  ( .A1(
        CipherErrorVec[14]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n33 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n34 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U17  ( .A1(
        CipherErrorVec[12]), .A2(CipherErrorVec[13]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n32 ), .B(
        AddRoundKeyOutput[17]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n30 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U13  ( .A(
        AddRoundKeyOutput[16]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n28 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U12  ( .A1(
        CipherErrorVec[13]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n27 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U11  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U10  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n24 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n23 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n31 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n23 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U8  ( .A(
        AddRoundKeyOutput[19]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n22 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U7  ( .A1(
        CipherErrorVec[12]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n22 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U6  ( .A1(
        CipherErrorVec[13]), .A2(CipherErrorVec[14]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U5  ( .A(
        AddRoundKeyOutput[18]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n20 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U4  ( .A1(
        CipherErrorVec[13]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U3  ( .A1(
        CipherErrorVec[14]), .A2(CipherErrorVec[12]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n25 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U22  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n36 ), .ZN(
        Red_PermutationInput[13]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n36 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n33 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n34 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U18  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n30 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n37 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U17  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n29 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n28 ), .B(
        AddRoundKeyOutput[16]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n31 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n28 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U14  ( .A(
        AddRoundKeyOutput[18]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n25 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n35 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U13  ( .A1(
        CipherErrorVec[13]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n24 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U12  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n23 ), .A2(
        CipherErrorVec[14]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n32 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n22 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n30 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U10  ( .A(
        AddRoundKeyOutput[19]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n21 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n22 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U9  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n23 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n21 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U8  ( .A1(
        CipherErrorVec[13]), .A2(CipherErrorVec[14]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n27 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U7  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n20 ), .B(
        AddRoundKeyOutput[17]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n32 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U6  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n19 ), .A2(
        CipherErrorVec[14]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U5  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n23 ), .A2(
        CipherErrorVec[13]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n19 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U4  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U3  ( .A(
        CipherErrorVec[12]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n36 ), .ZN(
        Red_PermutationInput[14]) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n36 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U19  ( .A(
        AddRoundKeyOutput[17]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n33 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n34 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U18  ( .A1(
        CipherErrorVec[14]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n33 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U17  ( .A1(
        CipherErrorVec[12]), .A2(CipherErrorVec[13]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U16  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n31 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n37 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U13  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n26 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U12  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n25 ), .B(
        AddRoundKeyOutput[18]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n28 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n24 ), .A2(
        CipherErrorVec[13]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U10  ( .A1(
        CipherErrorVec[12]), .A2(CipherErrorVec[14]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n24 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n29 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n30 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n27 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U8  ( .A(
        AddRoundKeyOutput[16]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n23 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n30 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U7  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n22 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U6  ( .A(
        CipherErrorVec[12]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n22 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U5  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n20 ), .B(
        AddRoundKeyOutput[19]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U4  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n21 ), .A2(
        CipherErrorVec[12]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U3  ( .A1(
        CipherErrorVec[13]), .A2(CipherErrorVec[14]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n35 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n34 ), .ZN(
        Red_PermutationInput[15]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U18  ( .A1(
        CipherErrorVec[17]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n33 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n34 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U17  ( .A1(
        CipherErrorVec[15]), .A2(CipherErrorVec[16]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n32 ), .B(
        AddRoundKeyOutput[21]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n30 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U13  ( .A(
        AddRoundKeyOutput[20]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n28 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U12  ( .A1(
        CipherErrorVec[16]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n27 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U11  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U10  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n24 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n23 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n31 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n23 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U8  ( .A(
        AddRoundKeyOutput[23]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n22 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U7  ( .A1(
        CipherErrorVec[15]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n22 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U6  ( .A1(
        CipherErrorVec[16]), .A2(CipherErrorVec[17]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U5  ( .A(
        AddRoundKeyOutput[22]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n20 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U4  ( .A1(
        CipherErrorVec[16]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U3  ( .A1(
        CipherErrorVec[17]), .A2(CipherErrorVec[15]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n25 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U22  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n36 ), .ZN(
        Red_PermutationInput[16]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n36 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n33 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n34 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U18  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n30 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n37 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U17  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n29 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n28 ), .B(
        AddRoundKeyOutput[20]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n31 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n28 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U14  ( .A(
        AddRoundKeyOutput[22]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n25 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n35 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U13  ( .A1(
        CipherErrorVec[16]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n24 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U12  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n23 ), .A2(
        CipherErrorVec[17]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n32 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n22 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n30 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U10  ( .A(
        AddRoundKeyOutput[23]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n21 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n22 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U9  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n23 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n21 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U8  ( .A1(
        CipherErrorVec[16]), .A2(CipherErrorVec[17]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n27 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U7  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n20 ), .B(
        AddRoundKeyOutput[21]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n32 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U6  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n19 ), .A2(
        CipherErrorVec[17]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U5  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n23 ), .A2(
        CipherErrorVec[16]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n19 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U4  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U3  ( .A(
        CipherErrorVec[15]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n36 ), .ZN(
        Red_PermutationInput[17]) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n36 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U19  ( .A(
        AddRoundKeyOutput[21]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n33 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n34 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U18  ( .A1(
        CipherErrorVec[17]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n33 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U17  ( .A1(
        CipherErrorVec[15]), .A2(CipherErrorVec[16]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U16  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n31 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n37 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U13  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n26 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U12  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n25 ), .B(
        AddRoundKeyOutput[22]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n28 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n24 ), .A2(
        CipherErrorVec[16]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U10  ( .A1(
        CipherErrorVec[15]), .A2(CipherErrorVec[17]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n24 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n29 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n30 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n27 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U8  ( .A(
        AddRoundKeyOutput[20]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n23 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n30 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U7  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n22 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U6  ( .A(
        CipherErrorVec[15]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n22 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U5  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n20 ), .B(
        AddRoundKeyOutput[23]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U4  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n21 ), .A2(
        CipherErrorVec[15]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U3  ( .A1(
        CipherErrorVec[16]), .A2(CipherErrorVec[17]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n35 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n34 ), .ZN(
        Red_PermutationInput[18]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U18  ( .A1(
        CipherErrorVec[20]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n33 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n34 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U17  ( .A1(
        CipherErrorVec[18]), .A2(CipherErrorVec[19]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n32 ), .B(
        AddRoundKeyOutput[25]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n30 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U13  ( .A(
        AddRoundKeyOutput[24]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n28 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U12  ( .A1(
        CipherErrorVec[19]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n27 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U11  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U10  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n24 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n23 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n31 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n23 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U8  ( .A(
        AddRoundKeyOutput[27]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n22 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U7  ( .A1(
        CipherErrorVec[18]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n22 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U6  ( .A1(
        CipherErrorVec[19]), .A2(CipherErrorVec[20]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U5  ( .A(
        AddRoundKeyOutput[26]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n20 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U4  ( .A1(
        CipherErrorVec[19]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U3  ( .A1(
        CipherErrorVec[20]), .A2(CipherErrorVec[18]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n25 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U22  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n36 ), .ZN(
        Red_PermutationInput[19]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n36 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n33 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n34 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U18  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n30 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n37 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U17  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n29 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n28 ), .B(
        AddRoundKeyOutput[24]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n31 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n28 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U14  ( .A(
        AddRoundKeyOutput[26]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n25 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n35 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U13  ( .A1(
        CipherErrorVec[19]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n24 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U12  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n23 ), .A2(
        CipherErrorVec[20]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n32 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n22 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n30 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U10  ( .A(
        AddRoundKeyOutput[27]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n21 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n22 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U9  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n23 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n21 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U8  ( .A1(
        CipherErrorVec[19]), .A2(CipherErrorVec[20]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n27 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U7  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n20 ), .B(
        AddRoundKeyOutput[25]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n32 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U6  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n19 ), .A2(
        CipherErrorVec[20]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U5  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n23 ), .A2(
        CipherErrorVec[19]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n19 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U4  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U3  ( .A(
        CipherErrorVec[18]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n36 ), .ZN(
        Red_PermutationInput[20]) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n36 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U19  ( .A(
        AddRoundKeyOutput[25]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n33 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n34 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U18  ( .A1(
        CipherErrorVec[20]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n33 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U17  ( .A1(
        CipherErrorVec[18]), .A2(CipherErrorVec[19]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U16  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n31 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n37 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U13  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n26 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U12  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n25 ), .B(
        AddRoundKeyOutput[26]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n28 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n24 ), .A2(
        CipherErrorVec[19]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U10  ( .A1(
        CipherErrorVec[18]), .A2(CipherErrorVec[20]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n24 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n29 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n30 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n27 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U8  ( .A(
        AddRoundKeyOutput[24]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n23 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n30 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U7  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n22 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U6  ( .A(
        CipherErrorVec[18]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n22 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U5  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n20 ), .B(
        AddRoundKeyOutput[27]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U4  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n21 ), .A2(
        CipherErrorVec[18]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U3  ( .A1(
        CipherErrorVec[19]), .A2(CipherErrorVec[20]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n35 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n34 ), .ZN(
        Red_PermutationInput[21]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U18  ( .A1(
        CipherErrorVec[23]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n33 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n34 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U17  ( .A1(
        CipherErrorVec[21]), .A2(CipherErrorVec[22]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n32 ), .B(
        AddRoundKeyOutput[29]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n30 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U13  ( .A(
        AddRoundKeyOutput[28]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n28 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U12  ( .A1(
        CipherErrorVec[22]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n27 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U11  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U10  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n24 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n23 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n31 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n23 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U8  ( .A(
        AddRoundKeyOutput[31]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n22 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U7  ( .A1(
        CipherErrorVec[21]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n22 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U6  ( .A1(
        CipherErrorVec[22]), .A2(CipherErrorVec[23]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U5  ( .A(
        AddRoundKeyOutput[30]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n20 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U4  ( .A1(
        CipherErrorVec[22]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U3  ( .A1(
        CipherErrorVec[23]), .A2(CipherErrorVec[21]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n25 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U22  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n36 ), .ZN(
        Red_PermutationInput[22]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n36 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n33 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n34 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U18  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n30 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n37 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U17  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n29 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n28 ), .B(
        AddRoundKeyOutput[28]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n31 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n28 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U14  ( .A(
        AddRoundKeyOutput[30]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n25 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n35 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U13  ( .A1(
        CipherErrorVec[22]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n24 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U12  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n23 ), .A2(
        CipherErrorVec[23]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n32 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n22 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n30 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U10  ( .A(
        AddRoundKeyOutput[31]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n21 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n22 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U9  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n23 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n21 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U8  ( .A1(
        CipherErrorVec[22]), .A2(CipherErrorVec[23]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n27 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U7  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n20 ), .B(
        AddRoundKeyOutput[29]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n32 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U6  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n19 ), .A2(
        CipherErrorVec[23]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U5  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n23 ), .A2(
        CipherErrorVec[22]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n19 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U4  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U3  ( .A(
        CipherErrorVec[21]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n36 ), .ZN(
        Red_PermutationInput[23]) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n36 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U19  ( .A(
        AddRoundKeyOutput[29]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n33 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n34 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U18  ( .A1(
        CipherErrorVec[23]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n33 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U17  ( .A1(
        CipherErrorVec[21]), .A2(CipherErrorVec[22]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U16  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n31 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n37 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U13  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n26 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U12  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n25 ), .B(
        AddRoundKeyOutput[30]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n28 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n24 ), .A2(
        CipherErrorVec[22]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U10  ( .A1(
        CipherErrorVec[21]), .A2(CipherErrorVec[23]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n24 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n29 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n30 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n27 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U8  ( .A(
        AddRoundKeyOutput[28]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n23 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n30 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U7  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n22 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U6  ( .A(
        CipherErrorVec[21]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n22 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U5  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n20 ), .B(
        AddRoundKeyOutput[31]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U4  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n21 ), .A2(
        CipherErrorVec[21]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U3  ( .A1(
        CipherErrorVec[22]), .A2(CipherErrorVec[23]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n35 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n34 ), .ZN(
        Red_PermutationInput[24]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U18  ( .A1(
        CipherErrorVec[26]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n33 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n34 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U17  ( .A1(
        CipherErrorVec[24]), .A2(CipherErrorVec[25]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n32 ), .B(
        AddRoundKeyOutput[33]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n30 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U13  ( .A(
        AddRoundKeyOutput[32]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n28 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U12  ( .A1(
        CipherErrorVec[25]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n27 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U11  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U10  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n24 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n23 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n31 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n23 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U8  ( .A(
        AddRoundKeyOutput[35]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n22 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U7  ( .A1(
        CipherErrorVec[24]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n22 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U6  ( .A1(
        CipherErrorVec[25]), .A2(CipherErrorVec[26]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U5  ( .A(
        AddRoundKeyOutput[34]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n20 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U4  ( .A1(
        CipherErrorVec[25]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U3  ( .A1(
        CipherErrorVec[26]), .A2(CipherErrorVec[24]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n25 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U22  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n36 ), .ZN(
        Red_PermutationInput[25]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n36 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n33 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n34 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U18  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n30 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n37 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U17  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n29 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n28 ), .B(
        AddRoundKeyOutput[32]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n31 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n28 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U14  ( .A(
        AddRoundKeyOutput[34]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n25 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n35 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U13  ( .A1(
        CipherErrorVec[25]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n24 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U12  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n23 ), .A2(
        CipherErrorVec[26]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n32 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n22 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n30 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U10  ( .A(
        AddRoundKeyOutput[35]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n21 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n22 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U9  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n23 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n21 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U8  ( .A1(
        CipherErrorVec[25]), .A2(CipherErrorVec[26]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n27 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U7  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n20 ), .B(
        AddRoundKeyOutput[33]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n32 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U6  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n19 ), .A2(
        CipherErrorVec[26]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U5  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n23 ), .A2(
        CipherErrorVec[25]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n19 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U4  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U3  ( .A(
        CipherErrorVec[24]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n36 ), .ZN(
        Red_PermutationInput[26]) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n36 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U19  ( .A(
        AddRoundKeyOutput[33]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n33 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n34 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U18  ( .A1(
        CipherErrorVec[26]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n33 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U17  ( .A1(
        CipherErrorVec[24]), .A2(CipherErrorVec[25]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U16  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n31 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n37 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U13  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n26 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U12  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n25 ), .B(
        AddRoundKeyOutput[34]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n28 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n24 ), .A2(
        CipherErrorVec[25]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U10  ( .A1(
        CipherErrorVec[24]), .A2(CipherErrorVec[26]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n24 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n29 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n30 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n27 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U8  ( .A(
        AddRoundKeyOutput[32]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n23 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n30 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U7  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n22 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U6  ( .A(
        CipherErrorVec[24]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n22 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U5  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n20 ), .B(
        AddRoundKeyOutput[35]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U4  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n21 ), .A2(
        CipherErrorVec[24]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U3  ( .A1(
        CipherErrorVec[25]), .A2(CipherErrorVec[26]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n35 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n34 ), .ZN(
        Red_PermutationInput[27]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U18  ( .A1(
        CipherErrorVec[29]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n33 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n34 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U17  ( .A1(
        CipherErrorVec[27]), .A2(CipherErrorVec[28]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n32 ), .B(
        AddRoundKeyOutput[37]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n30 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U13  ( .A(
        AddRoundKeyOutput[36]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n28 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U12  ( .A1(
        CipherErrorVec[28]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n27 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U11  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U10  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n24 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n23 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n31 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n23 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U8  ( .A(
        AddRoundKeyOutput[39]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n22 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U7  ( .A1(
        CipherErrorVec[27]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n22 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U6  ( .A1(
        CipherErrorVec[28]), .A2(CipherErrorVec[29]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U5  ( .A(
        AddRoundKeyOutput[38]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n20 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U4  ( .A1(
        CipherErrorVec[28]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U3  ( .A1(
        CipherErrorVec[29]), .A2(CipherErrorVec[27]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n25 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U22  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n36 ), .ZN(
        Red_PermutationInput[28]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n36 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n33 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n34 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U18  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n30 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n37 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U17  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n29 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n28 ), .B(
        AddRoundKeyOutput[36]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n31 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n28 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U14  ( .A(
        AddRoundKeyOutput[38]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n25 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n35 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U13  ( .A1(
        CipherErrorVec[28]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n24 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U12  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n23 ), .A2(
        CipherErrorVec[29]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n32 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n22 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n30 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U10  ( .A(
        AddRoundKeyOutput[39]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n21 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n22 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U9  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n23 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n21 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U8  ( .A1(
        CipherErrorVec[28]), .A2(CipherErrorVec[29]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n27 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U7  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n20 ), .B(
        AddRoundKeyOutput[37]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n32 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U6  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n19 ), .A2(
        CipherErrorVec[29]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U5  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n23 ), .A2(
        CipherErrorVec[28]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n19 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U4  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U3  ( .A(
        CipherErrorVec[27]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n36 ), .ZN(
        Red_PermutationInput[29]) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n36 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U19  ( .A(
        AddRoundKeyOutput[37]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n33 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n34 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U18  ( .A1(
        CipherErrorVec[29]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n33 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U17  ( .A1(
        CipherErrorVec[27]), .A2(CipherErrorVec[28]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U16  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n31 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n37 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U13  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n26 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U12  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n25 ), .B(
        AddRoundKeyOutput[38]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n28 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n24 ), .A2(
        CipherErrorVec[28]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U10  ( .A1(
        CipherErrorVec[27]), .A2(CipherErrorVec[29]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n24 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n29 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n30 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n27 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U8  ( .A(
        AddRoundKeyOutput[36]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n23 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n30 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U7  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n22 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U6  ( .A(
        CipherErrorVec[27]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n22 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U5  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n20 ), .B(
        AddRoundKeyOutput[39]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U4  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n21 ), .A2(
        CipherErrorVec[27]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U3  ( .A1(
        CipherErrorVec[28]), .A2(CipherErrorVec[29]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n35 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n34 ), .ZN(
        Red_PermutationInput[30]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U18  ( .A1(
        CipherErrorVec[32]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n33 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n34 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U17  ( .A1(
        CipherErrorVec[30]), .A2(CipherErrorVec[31]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n32 ), .B(
        AddRoundKeyOutput[41]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n30 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U13  ( .A(
        AddRoundKeyOutput[40]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n28 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U12  ( .A1(
        CipherErrorVec[31]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n27 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U11  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U10  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n24 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n23 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n31 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n23 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U8  ( .A(
        AddRoundKeyOutput[43]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n22 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U7  ( .A1(
        CipherErrorVec[30]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n22 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U6  ( .A1(
        CipherErrorVec[31]), .A2(CipherErrorVec[32]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U5  ( .A(
        AddRoundKeyOutput[42]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n20 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U4  ( .A1(
        CipherErrorVec[31]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U3  ( .A1(
        CipherErrorVec[32]), .A2(CipherErrorVec[30]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n25 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U22  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n36 ), .ZN(
        Red_PermutationInput[31]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n36 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n33 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n34 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U18  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n30 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n37 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U17  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n29 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n28 ), .B(
        AddRoundKeyOutput[40]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n31 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n28 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U14  ( .A(
        AddRoundKeyOutput[42]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n25 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n35 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U13  ( .A1(
        CipherErrorVec[31]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n24 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U12  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n23 ), .A2(
        CipherErrorVec[32]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n32 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n22 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n30 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U10  ( .A(
        AddRoundKeyOutput[43]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n21 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n22 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U9  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n23 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n21 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U8  ( .A1(
        CipherErrorVec[31]), .A2(CipherErrorVec[32]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n27 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U7  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n20 ), .B(
        AddRoundKeyOutput[41]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n32 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U6  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n19 ), .A2(
        CipherErrorVec[32]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U5  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n23 ), .A2(
        CipherErrorVec[31]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n19 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U4  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U3  ( .A(
        CipherErrorVec[30]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n36 ), .ZN(
        Red_PermutationInput[32]) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n36 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U19  ( .A(
        AddRoundKeyOutput[41]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n33 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n34 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U18  ( .A1(
        CipherErrorVec[32]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n33 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U17  ( .A1(
        CipherErrorVec[30]), .A2(CipherErrorVec[31]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U16  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n31 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n37 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U13  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n26 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U12  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n25 ), .B(
        AddRoundKeyOutput[42]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n28 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n24 ), .A2(
        CipherErrorVec[31]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U10  ( .A1(
        CipherErrorVec[30]), .A2(CipherErrorVec[32]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n24 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n29 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n30 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n27 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U8  ( .A(
        AddRoundKeyOutput[40]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n23 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n30 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U7  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n22 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U6  ( .A(
        CipherErrorVec[30]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n22 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U5  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n20 ), .B(
        AddRoundKeyOutput[43]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U4  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n21 ), .A2(
        CipherErrorVec[30]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U3  ( .A1(
        CipherErrorVec[31]), .A2(CipherErrorVec[32]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n35 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n34 ), .ZN(
        Red_PermutationInput[33]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U18  ( .A1(
        CipherErrorVec[35]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n33 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n34 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U17  ( .A1(
        CipherErrorVec[33]), .A2(CipherErrorVec[34]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n32 ), .B(
        AddRoundKeyOutput[45]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n30 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U13  ( .A(
        AddRoundKeyOutput[44]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n28 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U12  ( .A1(
        CipherErrorVec[34]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n27 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U11  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U10  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n24 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n23 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n31 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n23 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U8  ( .A(
        AddRoundKeyOutput[47]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n22 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U7  ( .A1(
        CipherErrorVec[33]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n22 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U6  ( .A1(
        CipherErrorVec[34]), .A2(CipherErrorVec[35]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U5  ( .A(
        AddRoundKeyOutput[46]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n20 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U4  ( .A1(
        CipherErrorVec[34]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U3  ( .A1(
        CipherErrorVec[35]), .A2(CipherErrorVec[33]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n25 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U22  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n36 ), .ZN(
        Red_PermutationInput[34]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n36 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n33 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n34 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U18  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n30 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n37 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U17  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n29 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n28 ), .B(
        AddRoundKeyOutput[44]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n31 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n28 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U14  ( .A(
        AddRoundKeyOutput[46]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n25 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n35 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U13  ( .A1(
        CipherErrorVec[34]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n24 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U12  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n23 ), .A2(
        CipherErrorVec[35]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n32 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n22 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n30 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U10  ( .A(
        AddRoundKeyOutput[47]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n21 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n22 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U9  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n23 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n21 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U8  ( .A1(
        CipherErrorVec[34]), .A2(CipherErrorVec[35]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n27 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U7  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n20 ), .B(
        AddRoundKeyOutput[45]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n32 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U6  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n19 ), .A2(
        CipherErrorVec[35]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U5  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n23 ), .A2(
        CipherErrorVec[34]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n19 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U4  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U3  ( .A(
        CipherErrorVec[33]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n36 ), .ZN(
        Red_PermutationInput[35]) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n36 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U19  ( .A(
        AddRoundKeyOutput[45]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n33 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n34 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U18  ( .A1(
        CipherErrorVec[35]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n33 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U17  ( .A1(
        CipherErrorVec[33]), .A2(CipherErrorVec[34]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U16  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n31 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n37 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U13  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n26 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U12  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n25 ), .B(
        AddRoundKeyOutput[46]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n28 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n24 ), .A2(
        CipherErrorVec[34]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U10  ( .A1(
        CipherErrorVec[33]), .A2(CipherErrorVec[35]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n24 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n29 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n30 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n27 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U8  ( .A(
        AddRoundKeyOutput[44]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n23 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n30 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U7  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n22 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U6  ( .A(
        CipherErrorVec[33]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n22 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U5  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n20 ), .B(
        AddRoundKeyOutput[47]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U4  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n21 ), .A2(
        CipherErrorVec[33]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U3  ( .A1(
        CipherErrorVec[34]), .A2(CipherErrorVec[35]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n35 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n34 ), .ZN(
        Red_PermutationInput[36]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U18  ( .A1(
        CipherErrorVec[38]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n33 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n34 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U17  ( .A1(
        CipherErrorVec[36]), .A2(CipherErrorVec[37]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n32 ), .B(
        AddRoundKeyOutput[49]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n30 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U13  ( .A(
        AddRoundKeyOutput[48]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n28 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U12  ( .A1(
        CipherErrorVec[37]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n27 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U11  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U10  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n24 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n23 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n31 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n23 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U8  ( .A(
        AddRoundKeyOutput[51]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n22 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U7  ( .A1(
        CipherErrorVec[36]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n22 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U6  ( .A1(
        CipherErrorVec[37]), .A2(CipherErrorVec[38]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U5  ( .A(
        AddRoundKeyOutput[50]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n20 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U4  ( .A1(
        CipherErrorVec[37]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U3  ( .A1(
        CipherErrorVec[38]), .A2(CipherErrorVec[36]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n25 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U22  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n36 ), .ZN(
        Red_PermutationInput[37]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n36 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n33 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n34 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U18  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n30 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n37 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U17  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n29 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n28 ), .B(
        AddRoundKeyOutput[48]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n31 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n28 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U14  ( .A(
        AddRoundKeyOutput[50]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n25 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n35 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U13  ( .A1(
        CipherErrorVec[37]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n24 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U12  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n23 ), .A2(
        CipherErrorVec[38]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n32 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n22 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n30 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U10  ( .A(
        AddRoundKeyOutput[51]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n21 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n22 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U9  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n23 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n21 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U8  ( .A1(
        CipherErrorVec[37]), .A2(CipherErrorVec[38]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n27 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U7  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n20 ), .B(
        AddRoundKeyOutput[49]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n32 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U6  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n19 ), .A2(
        CipherErrorVec[38]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U5  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n23 ), .A2(
        CipherErrorVec[37]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n19 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U4  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U3  ( .A(
        CipherErrorVec[36]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n36 ), .ZN(
        Red_PermutationInput[38]) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n36 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U19  ( .A(
        AddRoundKeyOutput[49]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n33 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n34 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U18  ( .A1(
        CipherErrorVec[38]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n33 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U17  ( .A1(
        CipherErrorVec[36]), .A2(CipherErrorVec[37]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U16  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n31 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n37 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U13  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n26 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U12  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n25 ), .B(
        AddRoundKeyOutput[50]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n28 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n24 ), .A2(
        CipherErrorVec[37]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U10  ( .A1(
        CipherErrorVec[36]), .A2(CipherErrorVec[38]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n24 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n29 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n30 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n27 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U8  ( .A(
        AddRoundKeyOutput[48]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n23 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n30 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U7  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n22 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U6  ( .A(
        CipherErrorVec[36]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n22 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U5  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n20 ), .B(
        AddRoundKeyOutput[51]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U4  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n21 ), .A2(
        CipherErrorVec[36]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U3  ( .A1(
        CipherErrorVec[37]), .A2(CipherErrorVec[38]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n35 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n34 ), .ZN(
        Red_PermutationInput[39]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U18  ( .A1(
        CipherErrorVec[41]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n33 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n34 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U17  ( .A1(
        CipherErrorVec[39]), .A2(CipherErrorVec[40]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n32 ), .B(
        AddRoundKeyOutput[53]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n30 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U13  ( .A(
        AddRoundKeyOutput[52]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n28 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U12  ( .A1(
        CipherErrorVec[40]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n27 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U11  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U10  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n24 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n23 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n31 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n23 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U8  ( .A(
        AddRoundKeyOutput[55]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n22 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U7  ( .A1(
        CipherErrorVec[39]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n22 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U6  ( .A1(
        CipherErrorVec[40]), .A2(CipherErrorVec[41]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U5  ( .A(
        AddRoundKeyOutput[54]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n20 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U4  ( .A1(
        CipherErrorVec[40]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U3  ( .A1(
        CipherErrorVec[41]), .A2(CipherErrorVec[39]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n25 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U22  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n36 ), .ZN(
        Red_PermutationInput[40]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n36 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n33 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n34 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U18  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n30 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n37 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U17  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n29 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n28 ), .B(
        AddRoundKeyOutput[52]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n31 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n28 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U14  ( .A(
        AddRoundKeyOutput[54]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n25 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n35 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U13  ( .A1(
        CipherErrorVec[40]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n24 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U12  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n23 ), .A2(
        CipherErrorVec[41]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n32 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n22 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n30 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U10  ( .A(
        AddRoundKeyOutput[55]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n21 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n22 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U9  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n23 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n21 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U8  ( .A1(
        CipherErrorVec[40]), .A2(CipherErrorVec[41]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n27 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U7  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n20 ), .B(
        AddRoundKeyOutput[53]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n32 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U6  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n19 ), .A2(
        CipherErrorVec[41]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U5  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n23 ), .A2(
        CipherErrorVec[40]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n19 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U4  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U3  ( .A(
        CipherErrorVec[39]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n36 ), .ZN(
        Red_PermutationInput[41]) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n36 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U19  ( .A(
        AddRoundKeyOutput[53]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n33 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n34 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U18  ( .A1(
        CipherErrorVec[41]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n33 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U17  ( .A1(
        CipherErrorVec[39]), .A2(CipherErrorVec[40]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U16  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n31 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n37 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U13  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n26 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U12  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n25 ), .B(
        AddRoundKeyOutput[54]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n28 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n24 ), .A2(
        CipherErrorVec[40]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U10  ( .A1(
        CipherErrorVec[39]), .A2(CipherErrorVec[41]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n24 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n29 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n30 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n27 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U8  ( .A(
        AddRoundKeyOutput[52]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n23 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n30 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U7  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n22 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U6  ( .A(
        CipherErrorVec[39]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n22 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U5  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n20 ), .B(
        AddRoundKeyOutput[55]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U4  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n21 ), .A2(
        CipherErrorVec[39]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U3  ( .A1(
        CipherErrorVec[40]), .A2(CipherErrorVec[41]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n35 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n34 ), .ZN(
        Red_PermutationInput[42]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U18  ( .A1(
        CipherErrorVec[44]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n33 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n34 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U17  ( .A1(
        CipherErrorVec[42]), .A2(CipherErrorVec[43]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n32 ), .B(
        AddRoundKeyOutput[57]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n30 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U13  ( .A(
        AddRoundKeyOutput[56]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n28 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U12  ( .A1(
        CipherErrorVec[43]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n27 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U11  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U10  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n24 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n23 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n31 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n23 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U8  ( .A(
        AddRoundKeyOutput[59]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n22 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U7  ( .A1(
        CipherErrorVec[42]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n22 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U6  ( .A1(
        CipherErrorVec[43]), .A2(CipherErrorVec[44]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U5  ( .A(
        AddRoundKeyOutput[58]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n20 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U4  ( .A1(
        CipherErrorVec[43]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U3  ( .A1(
        CipherErrorVec[44]), .A2(CipherErrorVec[42]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n25 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U22  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n36 ), .ZN(
        Red_PermutationInput[43]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n36 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n33 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n34 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U18  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n30 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n37 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U17  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n29 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n28 ), .B(
        AddRoundKeyOutput[56]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n31 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n28 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U14  ( .A(
        AddRoundKeyOutput[58]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n25 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n35 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U13  ( .A1(
        CipherErrorVec[43]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n24 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U12  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n23 ), .A2(
        CipherErrorVec[44]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n32 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n22 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n30 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U10  ( .A(
        AddRoundKeyOutput[59]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n21 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n22 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U9  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n23 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n21 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U8  ( .A1(
        CipherErrorVec[43]), .A2(CipherErrorVec[44]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n27 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U7  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n20 ), .B(
        AddRoundKeyOutput[57]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n32 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U6  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n19 ), .A2(
        CipherErrorVec[44]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U5  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n23 ), .A2(
        CipherErrorVec[43]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n19 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U4  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U3  ( .A(
        CipherErrorVec[42]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n36 ), .ZN(
        Red_PermutationInput[44]) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n36 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U19  ( .A(
        AddRoundKeyOutput[57]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n33 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n34 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U18  ( .A1(
        CipherErrorVec[44]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n33 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U17  ( .A1(
        CipherErrorVec[42]), .A2(CipherErrorVec[43]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U16  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n31 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n37 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U13  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n26 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U12  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n25 ), .B(
        AddRoundKeyOutput[58]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n28 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n24 ), .A2(
        CipherErrorVec[43]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U10  ( .A1(
        CipherErrorVec[42]), .A2(CipherErrorVec[44]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n24 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n29 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n30 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n27 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U8  ( .A(
        AddRoundKeyOutput[56]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n23 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n30 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U7  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n22 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U6  ( .A(
        CipherErrorVec[42]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n22 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U5  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n20 ), .B(
        AddRoundKeyOutput[59]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U4  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n21 ), .A2(
        CipherErrorVec[42]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U3  ( .A1(
        CipherErrorVec[43]), .A2(CipherErrorVec[44]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n35 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n34 ), .ZN(
        Red_PermutationInput[45]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U18  ( .A1(
        CipherErrorVec[47]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n33 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n34 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U17  ( .A1(
        CipherErrorVec[45]), .A2(CipherErrorVec[46]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n32 ), .B(
        AddRoundKeyOutput[61]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n30 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U13  ( .A(
        AddRoundKeyOutput[60]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n28 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U12  ( .A1(
        CipherErrorVec[46]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n27 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U11  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U10  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n24 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n23 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n31 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n23 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U8  ( .A(
        AddRoundKeyOutput[63]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n22 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U7  ( .A1(
        CipherErrorVec[45]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n22 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U6  ( .A1(
        CipherErrorVec[46]), .A2(CipherErrorVec[47]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n21 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U5  ( .A(
        AddRoundKeyOutput[62]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n20 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U4  ( .A1(
        CipherErrorVec[46]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n25 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U3  ( .A1(
        CipherErrorVec[47]), .A2(CipherErrorVec[45]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n25 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U22  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n36 ), .ZN(
        Red_PermutationInput[46]) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n36 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n33 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n34 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U19  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n33 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U18  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n30 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n29 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n37 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U17  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n31 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n29 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U16  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n28 ), .B(
        AddRoundKeyOutput[60]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n31 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n28 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U14  ( .A(
        AddRoundKeyOutput[62]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n25 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n35 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U13  ( .A1(
        CipherErrorVec[46]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n24 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U12  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n23 ), .A2(
        CipherErrorVec[47]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n24 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n32 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n22 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n30 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U10  ( .A(
        AddRoundKeyOutput[63]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n21 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n22 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U9  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n23 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n27 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n21 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U8  ( .A1(
        CipherErrorVec[46]), .A2(CipherErrorVec[47]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n27 ) );
  XNOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U7  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n20 ), .B(
        AddRoundKeyOutput[61]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n32 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U6  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n19 ), .A2(
        CipherErrorVec[47]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U5  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n23 ), .A2(
        CipherErrorVec[46]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n19 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U4  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U3  ( .A(
        CipherErrorVec[45]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n26 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U21  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n37 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n36 ), .ZN(
        Red_PermutationInput[47]) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U20  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n35 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n34 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n36 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U19  ( .A(
        AddRoundKeyOutput[61]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n33 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n34 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U18  ( .A1(
        CipherErrorVec[47]), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n32 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n33 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U17  ( .A1(
        CipherErrorVec[45]), .A2(CipherErrorVec[46]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n32 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U16  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n31 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n30 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n35 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U15  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n29 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n31 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U14  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n27 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n26 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n37 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U13  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n28 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n26 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U12  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n25 ), .B(
        AddRoundKeyOutput[62]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n28 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U11  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n24 ), .A2(
        CipherErrorVec[46]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n25 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U10  ( .A1(
        CipherErrorVec[45]), .A2(CipherErrorVec[47]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n24 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U9  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n29 ), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n30 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n27 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U8  ( .A(
        AddRoundKeyOutput[60]), .B(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n23 ), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n30 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U7  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n22 ), .A2(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n21 ), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n23 ) );
  INV_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U6  ( .A(
        CipherErrorVec[45]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n22 ) );
  XOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U5  ( .A(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n20 ), .B(
        AddRoundKeyOutput[63]), .Z(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n29 ) );
  NOR2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U4  ( .A1(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n21 ), .A2(
        CipherErrorVec[45]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n20 ) );
  NAND2_X1 \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U3  ( .A1(
        CipherErrorVec[46]), .A2(CipherErrorVec[47]), .ZN(
        \SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n21 ) );
  DFF_X1 \Red_StateReg_s_current_state_reg[0]  ( .D(Red_PermutationInput[0]), 
        .CK(clk), .Q(Red_Feedback[45]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[1]  ( .D(Red_PermutationInput[1]), 
        .CK(clk), .Q(Red_Feedback[46]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[2]  ( .D(Red_PermutationInput[2]), 
        .CK(clk), .Q(Red_Feedback[47]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[3]  ( .D(Red_PermutationInput[3]), 
        .CK(clk), .Q(Red_Feedback[36]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[4]  ( .D(Red_PermutationInput[4]), 
        .CK(clk), .Q(Red_Feedback[37]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[5]  ( .D(Red_PermutationInput[5]), 
        .CK(clk), .Q(Red_Feedback[38]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[6]  ( .D(Red_PermutationInput[6]), 
        .CK(clk), .Q(Red_Feedback[39]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[7]  ( .D(Red_PermutationInput[7]), 
        .CK(clk), .Q(Red_Feedback[40]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[8]  ( .D(Red_PermutationInput[8]), 
        .CK(clk), .Q(Red_Feedback[41]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[9]  ( .D(Red_PermutationInput[9]), 
        .CK(clk), .Q(Red_Feedback[42]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[10]  ( .D(Red_PermutationInput[10]), 
        .CK(clk), .Q(Red_Feedback[43]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[11]  ( .D(Red_PermutationInput[11]), 
        .CK(clk), .Q(Red_Feedback[44]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[12]  ( .D(Red_PermutationInput[12]), 
        .CK(clk), .Q(Red_Feedback[24]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[13]  ( .D(Red_PermutationInput[13]), 
        .CK(clk), .Q(Red_Feedback[25]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[14]  ( .D(Red_PermutationInput[14]), 
        .CK(clk), .Q(Red_Feedback[26]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[15]  ( .D(Red_PermutationInput[15]), 
        .CK(clk), .Q(Red_Feedback[33]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[16]  ( .D(Red_PermutationInput[16]), 
        .CK(clk), .Q(Red_Feedback[34]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[17]  ( .D(Red_PermutationInput[17]), 
        .CK(clk), .Q(Red_Feedback[35]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[18]  ( .D(Red_PermutationInput[18]), 
        .CK(clk), .Q(Red_Feedback[30]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[19]  ( .D(Red_PermutationInput[19]), 
        .CK(clk), .Q(Red_Feedback[31]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[20]  ( .D(Red_PermutationInput[20]), 
        .CK(clk), .Q(Red_Feedback[32]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[21]  ( .D(Red_PermutationInput[21]), 
        .CK(clk), .Q(Red_Feedback[27]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[22]  ( .D(Red_PermutationInput[22]), 
        .CK(clk), .Q(Red_Feedback[28]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[23]  ( .D(Red_PermutationInput[23]), 
        .CK(clk), .Q(Red_Feedback[29]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[24]  ( .D(Red_PermutationInput[24]), 
        .CK(clk), .Q(Red_Feedback[12]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[25]  ( .D(Red_PermutationInput[25]), 
        .CK(clk), .Q(Red_Feedback[13]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[26]  ( .D(Red_PermutationInput[26]), 
        .CK(clk), .Q(Red_Feedback[14]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[27]  ( .D(Red_PermutationInput[27]), 
        .CK(clk), .Q(Red_Feedback[21]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[28]  ( .D(Red_PermutationInput[28]), 
        .CK(clk), .Q(Red_Feedback[22]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[29]  ( .D(Red_PermutationInput[29]), 
        .CK(clk), .Q(Red_Feedback[23]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[30]  ( .D(Red_PermutationInput[30]), 
        .CK(clk), .Q(Red_Feedback[18]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[31]  ( .D(Red_PermutationInput[31]), 
        .CK(clk), .Q(Red_Feedback[19]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[32]  ( .D(Red_PermutationInput[32]), 
        .CK(clk), .Q(Red_Feedback[20]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[33]  ( .D(Red_PermutationInput[33]), 
        .CK(clk), .Q(Red_Feedback[15]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[34]  ( .D(Red_PermutationInput[34]), 
        .CK(clk), .Q(Red_Feedback[16]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[35]  ( .D(Red_PermutationInput[35]), 
        .CK(clk), .Q(Red_Feedback[17]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[36]  ( .D(Red_PermutationInput[36]), 
        .CK(clk), .Q(Red_Feedback[3]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[37]  ( .D(Red_PermutationInput[37]), 
        .CK(clk), .Q(Red_Feedback[4]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[38]  ( .D(Red_PermutationInput[38]), 
        .CK(clk), .Q(Red_Feedback[5]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[39]  ( .D(Red_PermutationInput[39]), 
        .CK(clk), .Q(Red_Feedback[6]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[40]  ( .D(Red_PermutationInput[40]), 
        .CK(clk), .Q(Red_Feedback[7]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[41]  ( .D(Red_PermutationInput[41]), 
        .CK(clk), .Q(Red_Feedback[8]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[42]  ( .D(Red_PermutationInput[42]), 
        .CK(clk), .Q(Red_Feedback[9]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[43]  ( .D(Red_PermutationInput[43]), 
        .CK(clk), .Q(Red_Feedback[10]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[44]  ( .D(Red_PermutationInput[44]), 
        .CK(clk), .Q(Red_Feedback[11]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[45]  ( .D(Red_PermutationInput[45]), 
        .CK(clk), .Q(Red_Feedback[0]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[46]  ( .D(Red_PermutationInput[46]), 
        .CK(clk), .Q(Red_Feedback[1]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[47]  ( .D(Red_PermutationInput[47]), 
        .CK(clk), .Q(Red_Feedback[2]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_0_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_0_LFInst_0_n2 ), .B(Feedback[1]), .ZN(
        FeedbackF[0]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_0_LFInst_0_U3  ( .A(Feedback[2]), .B(
        Feedback[0]), .ZN(\StateRegOutputF_inst2_LFInst_0_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_0_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_0_LFInst_1_n2 ), .B(Feedback[1]), .ZN(
        FeedbackF[1]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_0_LFInst_1_U3  ( .A(Feedback[3]), .B(
        Feedback[0]), .ZN(\StateRegOutputF_inst2_LFInst_0_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_0_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_0_LFInst_2_n2 ), .B(Feedback[2]), .ZN(
        FeedbackF[2]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_0_LFInst_2_U3  ( .A(Feedback[3]), .B(
        Feedback[0]), .ZN(\StateRegOutputF_inst2_LFInst_0_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_1_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_1_LFInst_0_n2 ), .B(Feedback[5]), .ZN(
        FeedbackF[3]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_1_LFInst_0_U3  ( .A(Feedback[6]), .B(
        Feedback[4]), .ZN(\StateRegOutputF_inst2_LFInst_1_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_1_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_1_LFInst_1_n2 ), .B(Feedback[5]), .ZN(
        FeedbackF[4]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_1_LFInst_1_U3  ( .A(Feedback[7]), .B(
        Feedback[4]), .ZN(\StateRegOutputF_inst2_LFInst_1_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_1_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_1_LFInst_2_n2 ), .B(Feedback[6]), .ZN(
        FeedbackF[5]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_1_LFInst_2_U3  ( .A(Feedback[7]), .B(
        Feedback[4]), .ZN(\StateRegOutputF_inst2_LFInst_1_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_2_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_2_LFInst_0_n2 ), .B(Feedback[9]), .ZN(
        FeedbackF[6]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_2_LFInst_0_U3  ( .A(Feedback[10]), 
        .B(Feedback[8]), .ZN(\StateRegOutputF_inst2_LFInst_2_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_2_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_2_LFInst_1_n2 ), .B(Feedback[9]), .ZN(
        FeedbackF[7]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_2_LFInst_1_U3  ( .A(Feedback[11]), 
        .B(Feedback[8]), .ZN(\StateRegOutputF_inst2_LFInst_2_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_2_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_2_LFInst_2_n2 ), .B(Feedback[10]), .ZN(
        FeedbackF[8]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_2_LFInst_2_U3  ( .A(Feedback[11]), 
        .B(Feedback[8]), .ZN(\StateRegOutputF_inst2_LFInst_2_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_3_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_3_LFInst_0_n2 ), .B(Feedback[13]), .ZN(
        FeedbackF[9]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_3_LFInst_0_U3  ( .A(Feedback[14]), 
        .B(Feedback[12]), .ZN(\StateRegOutputF_inst2_LFInst_3_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_3_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_3_LFInst_1_n2 ), .B(Feedback[13]), .ZN(
        FeedbackF[10]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_3_LFInst_1_U3  ( .A(Feedback[15]), 
        .B(Feedback[12]), .ZN(\StateRegOutputF_inst2_LFInst_3_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_3_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_3_LFInst_2_n2 ), .B(Feedback[14]), .ZN(
        FeedbackF[11]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_3_LFInst_2_U3  ( .A(Feedback[15]), 
        .B(Feedback[12]), .ZN(\StateRegOutputF_inst2_LFInst_3_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_4_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_4_LFInst_0_n2 ), .B(Feedback[17]), .ZN(
        FeedbackF[12]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_4_LFInst_0_U3  ( .A(Feedback[18]), 
        .B(Feedback[16]), .ZN(\StateRegOutputF_inst2_LFInst_4_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_4_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_4_LFInst_1_n2 ), .B(Feedback[17]), .ZN(
        FeedbackF[13]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_4_LFInst_1_U3  ( .A(Feedback[19]), 
        .B(Feedback[16]), .ZN(\StateRegOutputF_inst2_LFInst_4_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_4_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_4_LFInst_2_n2 ), .B(Feedback[18]), .ZN(
        FeedbackF[14]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_4_LFInst_2_U3  ( .A(Feedback[19]), 
        .B(Feedback[16]), .ZN(\StateRegOutputF_inst2_LFInst_4_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_5_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_5_LFInst_0_n2 ), .B(Feedback[21]), .ZN(
        FeedbackF[15]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_5_LFInst_0_U3  ( .A(Feedback[22]), 
        .B(Feedback[20]), .ZN(\StateRegOutputF_inst2_LFInst_5_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_5_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_5_LFInst_1_n2 ), .B(Feedback[21]), .ZN(
        FeedbackF[16]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_5_LFInst_1_U3  ( .A(Feedback[23]), 
        .B(Feedback[20]), .ZN(\StateRegOutputF_inst2_LFInst_5_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_5_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_5_LFInst_2_n2 ), .B(Feedback[22]), .ZN(
        FeedbackF[17]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_5_LFInst_2_U3  ( .A(Feedback[23]), 
        .B(Feedback[20]), .ZN(\StateRegOutputF_inst2_LFInst_5_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_6_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_6_LFInst_0_n2 ), .B(Feedback[25]), .ZN(
        FeedbackF[18]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_6_LFInst_0_U3  ( .A(Feedback[26]), 
        .B(Feedback[24]), .ZN(\StateRegOutputF_inst2_LFInst_6_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_6_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_6_LFInst_1_n2 ), .B(Feedback[25]), .ZN(
        FeedbackF[19]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_6_LFInst_1_U3  ( .A(Feedback[27]), 
        .B(Feedback[24]), .ZN(\StateRegOutputF_inst2_LFInst_6_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_6_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_6_LFInst_2_n2 ), .B(Feedback[26]), .ZN(
        FeedbackF[20]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_6_LFInst_2_U3  ( .A(Feedback[27]), 
        .B(Feedback[24]), .ZN(\StateRegOutputF_inst2_LFInst_6_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_7_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_7_LFInst_0_n2 ), .B(Feedback[29]), .ZN(
        FeedbackF[21]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_7_LFInst_0_U3  ( .A(Feedback[30]), 
        .B(Feedback[28]), .ZN(\StateRegOutputF_inst2_LFInst_7_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_7_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_7_LFInst_1_n2 ), .B(Feedback[29]), .ZN(
        FeedbackF[22]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_7_LFInst_1_U3  ( .A(Feedback[31]), 
        .B(Feedback[28]), .ZN(\StateRegOutputF_inst2_LFInst_7_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_7_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_7_LFInst_2_n2 ), .B(Feedback[30]), .ZN(
        FeedbackF[23]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_7_LFInst_2_U3  ( .A(Feedback[31]), 
        .B(Feedback[28]), .ZN(\StateRegOutputF_inst2_LFInst_7_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_8_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_8_LFInst_0_n2 ), .B(Feedback[33]), .ZN(
        FeedbackF[24]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_8_LFInst_0_U3  ( .A(Feedback[34]), 
        .B(Feedback[32]), .ZN(\StateRegOutputF_inst2_LFInst_8_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_8_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_8_LFInst_1_n2 ), .B(Feedback[33]), .ZN(
        FeedbackF[25]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_8_LFInst_1_U3  ( .A(Feedback[35]), 
        .B(Feedback[32]), .ZN(\StateRegOutputF_inst2_LFInst_8_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_8_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_8_LFInst_2_n2 ), .B(Feedback[34]), .ZN(
        FeedbackF[26]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_8_LFInst_2_U3  ( .A(Feedback[35]), 
        .B(Feedback[32]), .ZN(\StateRegOutputF_inst2_LFInst_8_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_9_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_9_LFInst_0_n2 ), .B(Feedback[37]), .ZN(
        FeedbackF[27]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_9_LFInst_0_U3  ( .A(Feedback[38]), 
        .B(Feedback[36]), .ZN(\StateRegOutputF_inst2_LFInst_9_LFInst_0_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_9_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_9_LFInst_1_n2 ), .B(Feedback[37]), .ZN(
        FeedbackF[28]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_9_LFInst_1_U3  ( .A(Feedback[39]), 
        .B(Feedback[36]), .ZN(\StateRegOutputF_inst2_LFInst_9_LFInst_1_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_9_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_9_LFInst_2_n2 ), .B(Feedback[38]), .ZN(
        FeedbackF[29]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_9_LFInst_2_U3  ( .A(Feedback[39]), 
        .B(Feedback[36]), .ZN(\StateRegOutputF_inst2_LFInst_9_LFInst_2_n2 ) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_10_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_10_LFInst_0_n2 ), .B(Feedback[41]), .ZN(
        FeedbackF[30]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_10_LFInst_0_U3  ( .A(Feedback[42]), 
        .B(Feedback[40]), .ZN(\StateRegOutputF_inst2_LFInst_10_LFInst_0_n2 )
         );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_10_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_10_LFInst_1_n2 ), .B(Feedback[41]), .ZN(
        FeedbackF[31]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_10_LFInst_1_U3  ( .A(Feedback[43]), 
        .B(Feedback[40]), .ZN(\StateRegOutputF_inst2_LFInst_10_LFInst_1_n2 )
         );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_10_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_10_LFInst_2_n2 ), .B(Feedback[42]), .ZN(
        FeedbackF[32]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_10_LFInst_2_U3  ( .A(Feedback[43]), 
        .B(Feedback[40]), .ZN(\StateRegOutputF_inst2_LFInst_10_LFInst_2_n2 )
         );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_11_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_11_LFInst_0_n2 ), .B(Feedback[45]), .ZN(
        FeedbackF[33]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_11_LFInst_0_U3  ( .A(Feedback[46]), 
        .B(Feedback[44]), .ZN(\StateRegOutputF_inst2_LFInst_11_LFInst_0_n2 )
         );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_11_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_11_LFInst_1_n2 ), .B(Feedback[45]), .ZN(
        FeedbackF[34]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_11_LFInst_1_U3  ( .A(Feedback[47]), 
        .B(Feedback[44]), .ZN(\StateRegOutputF_inst2_LFInst_11_LFInst_1_n2 )
         );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_11_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_11_LFInst_2_n2 ), .B(Feedback[46]), .ZN(
        FeedbackF[35]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_11_LFInst_2_U3  ( .A(Feedback[47]), 
        .B(Feedback[44]), .ZN(\StateRegOutputF_inst2_LFInst_11_LFInst_2_n2 )
         );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_12_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_12_LFInst_0_n2 ), .B(Feedback[49]), .ZN(
        FeedbackF[36]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_12_LFInst_0_U3  ( .A(Feedback[50]), 
        .B(Feedback[48]), .ZN(\StateRegOutputF_inst2_LFInst_12_LFInst_0_n2 )
         );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_12_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_12_LFInst_1_n2 ), .B(Feedback[49]), .ZN(
        FeedbackF[37]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_12_LFInst_1_U3  ( .A(Feedback[51]), 
        .B(Feedback[48]), .ZN(\StateRegOutputF_inst2_LFInst_12_LFInst_1_n2 )
         );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_12_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_12_LFInst_2_n2 ), .B(Feedback[50]), .ZN(
        FeedbackF[38]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_12_LFInst_2_U3  ( .A(Feedback[51]), 
        .B(Feedback[48]), .ZN(\StateRegOutputF_inst2_LFInst_12_LFInst_2_n2 )
         );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_13_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_13_LFInst_0_n2 ), .B(Feedback[53]), .ZN(
        FeedbackF[39]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_13_LFInst_0_U3  ( .A(Feedback[54]), 
        .B(Feedback[52]), .ZN(\StateRegOutputF_inst2_LFInst_13_LFInst_0_n2 )
         );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_13_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_13_LFInst_1_n2 ), .B(Feedback[53]), .ZN(
        FeedbackF[40]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_13_LFInst_1_U3  ( .A(Feedback[55]), 
        .B(Feedback[52]), .ZN(\StateRegOutputF_inst2_LFInst_13_LFInst_1_n2 )
         );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_13_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_13_LFInst_2_n2 ), .B(Feedback[54]), .ZN(
        FeedbackF[41]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_13_LFInst_2_U3  ( .A(Feedback[55]), 
        .B(Feedback[52]), .ZN(\StateRegOutputF_inst2_LFInst_13_LFInst_2_n2 )
         );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_14_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_14_LFInst_0_n2 ), .B(Feedback[57]), .ZN(
        FeedbackF[42]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_14_LFInst_0_U3  ( .A(Feedback[58]), 
        .B(Feedback[56]), .ZN(\StateRegOutputF_inst2_LFInst_14_LFInst_0_n2 )
         );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_14_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_14_LFInst_1_n2 ), .B(Feedback[57]), .ZN(
        FeedbackF[43]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_14_LFInst_1_U3  ( .A(Feedback[59]), 
        .B(Feedback[56]), .ZN(\StateRegOutputF_inst2_LFInst_14_LFInst_1_n2 )
         );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_14_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_14_LFInst_2_n2 ), .B(Feedback[58]), .ZN(
        FeedbackF[44]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_14_LFInst_2_U3  ( .A(Feedback[59]), 
        .B(Feedback[56]), .ZN(\StateRegOutputF_inst2_LFInst_14_LFInst_2_n2 )
         );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_15_LFInst_0_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_15_LFInst_0_n2 ), .B(Feedback[61]), .ZN(
        FeedbackF[45]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_15_LFInst_0_U3  ( .A(Feedback[62]), 
        .B(Feedback[60]), .ZN(\StateRegOutputF_inst2_LFInst_15_LFInst_0_n2 )
         );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_15_LFInst_1_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_15_LFInst_1_n2 ), .B(Feedback[61]), .ZN(
        FeedbackF[46]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_15_LFInst_1_U3  ( .A(Feedback[63]), 
        .B(Feedback[60]), .ZN(\StateRegOutputF_inst2_LFInst_15_LFInst_1_n2 )
         );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_15_LFInst_2_U4  ( .A(
        \StateRegOutputF_inst2_LFInst_15_LFInst_2_n2 ), .B(Feedback[62]), .ZN(
        FeedbackF[47]) );
  XNOR2_X1 \StateRegOutputF_inst2_LFInst_15_LFInst_2_U3  ( .A(Feedback[63]), 
        .B(Feedback[60]), .ZN(\StateRegOutputF_inst2_LFInst_15_LFInst_2_n2 )
         );
  XOR2_X1 \CipherErrorVecGen2_XORInst_0_0_U1  ( .A(FeedbackF[0]), .B(
        Red_Feedback[0]), .Z(CipherErrorVec2[0]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_0_1_U1  ( .A(FeedbackF[1]), .B(
        Red_Feedback[1]), .Z(CipherErrorVec2[1]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_0_2_U1  ( .A(FeedbackF[2]), .B(
        Red_Feedback[2]), .Z(CipherErrorVec2[2]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_1_0_U1  ( .A(FeedbackF[3]), .B(
        Red_Feedback[3]), .Z(CipherErrorVec2[3]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_1_1_U1  ( .A(FeedbackF[4]), .B(
        Red_Feedback[4]), .Z(CipherErrorVec2[4]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_1_2_U1  ( .A(FeedbackF[5]), .B(
        Red_Feedback[5]), .Z(CipherErrorVec2[5]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_2_0_U1  ( .A(FeedbackF[6]), .B(
        Red_Feedback[6]), .Z(CipherErrorVec2[6]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_2_1_U1  ( .A(FeedbackF[7]), .B(
        Red_Feedback[7]), .Z(CipherErrorVec2[7]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_2_2_U1  ( .A(FeedbackF[8]), .B(
        Red_Feedback[8]), .Z(CipherErrorVec2[8]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_3_0_U1  ( .A(FeedbackF[9]), .B(
        Red_Feedback[9]), .Z(CipherErrorVec2[9]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_3_1_U1  ( .A(FeedbackF[10]), .B(
        Red_Feedback[10]), .Z(CipherErrorVec2[10]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_3_2_U1  ( .A(FeedbackF[11]), .B(
        Red_Feedback[11]), .Z(CipherErrorVec2[11]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_4_0_U1  ( .A(FeedbackF[12]), .B(
        Red_Feedback[12]), .Z(CipherErrorVec2[12]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_4_1_U1  ( .A(FeedbackF[13]), .B(
        Red_Feedback[13]), .Z(CipherErrorVec2[13]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_4_2_U1  ( .A(FeedbackF[14]), .B(
        Red_Feedback[14]), .Z(CipherErrorVec2[14]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_5_0_U1  ( .A(FeedbackF[15]), .B(
        Red_Feedback[15]), .Z(CipherErrorVec2[15]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_5_1_U1  ( .A(FeedbackF[16]), .B(
        Red_Feedback[16]), .Z(CipherErrorVec2[16]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_5_2_U1  ( .A(FeedbackF[17]), .B(
        Red_Feedback[17]), .Z(CipherErrorVec2[17]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_6_0_U1  ( .A(FeedbackF[18]), .B(
        Red_Feedback[18]), .Z(CipherErrorVec2[18]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_6_1_U1  ( .A(FeedbackF[19]), .B(
        Red_Feedback[19]), .Z(CipherErrorVec2[19]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_6_2_U1  ( .A(FeedbackF[20]), .B(
        Red_Feedback[20]), .Z(CipherErrorVec2[20]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_7_0_U1  ( .A(FeedbackF[21]), .B(
        Red_Feedback[21]), .Z(CipherErrorVec2[21]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_7_1_U1  ( .A(FeedbackF[22]), .B(
        Red_Feedback[22]), .Z(CipherErrorVec2[22]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_7_2_U1  ( .A(FeedbackF[23]), .B(
        Red_Feedback[23]), .Z(CipherErrorVec2[23]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_8_0_U1  ( .A(FeedbackF[24]), .B(
        Red_Feedback[24]), .Z(CipherErrorVec2[24]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_8_1_U1  ( .A(FeedbackF[25]), .B(
        Red_Feedback[25]), .Z(CipherErrorVec2[25]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_8_2_U1  ( .A(FeedbackF[26]), .B(
        Red_Feedback[26]), .Z(CipherErrorVec2[26]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_9_0_U1  ( .A(FeedbackF[27]), .B(
        Red_Feedback[27]), .Z(CipherErrorVec2[27]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_9_1_U1  ( .A(FeedbackF[28]), .B(
        Red_Feedback[28]), .Z(CipherErrorVec2[28]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_9_2_U1  ( .A(FeedbackF[29]), .B(
        Red_Feedback[29]), .Z(CipherErrorVec2[29]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_10_0_U1  ( .A(FeedbackF[30]), .B(
        Red_Feedback[30]), .Z(CipherErrorVec2[30]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_10_1_U1  ( .A(FeedbackF[31]), .B(
        Red_Feedback[31]), .Z(CipherErrorVec2[31]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_10_2_U1  ( .A(FeedbackF[32]), .B(
        Red_Feedback[32]), .Z(CipherErrorVec2[32]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_11_0_U1  ( .A(FeedbackF[33]), .B(
        Red_Feedback[33]), .Z(CipherErrorVec2[33]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_11_1_U1  ( .A(FeedbackF[34]), .B(
        Red_Feedback[34]), .Z(CipherErrorVec2[34]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_11_2_U1  ( .A(FeedbackF[35]), .B(
        Red_Feedback[35]), .Z(CipherErrorVec2[35]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_12_0_U1  ( .A(FeedbackF[36]), .B(
        Red_Feedback[36]), .Z(CipherErrorVec2[36]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_12_1_U1  ( .A(FeedbackF[37]), .B(
        Red_Feedback[37]), .Z(CipherErrorVec2[37]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_12_2_U1  ( .A(FeedbackF[38]), .B(
        Red_Feedback[38]), .Z(CipherErrorVec2[38]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_13_0_U1  ( .A(FeedbackF[39]), .B(
        Red_Feedback[39]), .Z(CipherErrorVec2[39]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_13_1_U1  ( .A(FeedbackF[40]), .B(
        Red_Feedback[40]), .Z(CipherErrorVec2[40]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_13_2_U1  ( .A(FeedbackF[41]), .B(
        Red_Feedback[41]), .Z(CipherErrorVec2[41]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_14_0_U1  ( .A(FeedbackF[42]), .B(
        Red_Feedback[42]), .Z(CipherErrorVec2[42]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_14_1_U1  ( .A(FeedbackF[43]), .B(
        Red_Feedback[43]), .Z(CipherErrorVec2[43]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_14_2_U1  ( .A(FeedbackF[44]), .B(
        Red_Feedback[44]), .Z(CipherErrorVec2[44]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_15_0_U1  ( .A(FeedbackF[45]), .B(
        Red_Feedback[45]), .Z(CipherErrorVec2[45]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_15_1_U1  ( .A(FeedbackF[46]), .B(
        Red_Feedback[46]), .Z(CipherErrorVec2[46]) );
  XOR2_X1 \CipherErrorVecGen2_XORInst_15_2_U1  ( .A(FeedbackF[47]), .B(
        Red_Feedback[47]), .Z(CipherErrorVec2[47]) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U14  ( .A(Feedback[0]), 
        .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n27 ), .Z(Output[0])
         );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U13  ( .A1(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n26 ), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n27 ) );
  INV_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U12  ( .A(
        CipherErrorVec2[0]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U11  ( .A(Feedback[1]), 
        .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n24 ), .Z(Output[1])
         );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U10  ( .A1(
        CipherErrorVec2[2]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n23 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U9  ( .A1(
        CipherErrorVec2[1]), .A2(CipherErrorVec2[0]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n23 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U8  ( .A(Feedback[2]), 
        .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n22 ), .Z(Output[2])
         );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U7  ( .A1(
        CipherErrorVec2[1]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n22 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U6  ( .A1(
        CipherErrorVec2[2]), .A2(CipherErrorVec2[0]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n21 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U5  ( .A(Feedback[3]), 
        .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n20 ), .Z(Output[3])
         );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U4  ( .A1(
        CipherErrorVec2[0]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U3  ( .A1(
        CipherErrorVec2[2]), .A2(CipherErrorVec2[1]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n26 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U14  ( .A(Feedback[4]), 
        .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n27 ), .Z(Output[4])
         );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U13  ( .A1(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n26 ), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n27 ) );
  INV_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U12  ( .A(
        CipherErrorVec2[3]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U11  ( .A(Feedback[5]), 
        .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n24 ), .Z(Output[5])
         );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U10  ( .A1(
        CipherErrorVec2[5]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n23 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U9  ( .A1(
        CipherErrorVec2[4]), .A2(CipherErrorVec2[3]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n23 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U8  ( .A(Feedback[6]), 
        .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n22 ), .Z(Output[6])
         );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U7  ( .A1(
        CipherErrorVec2[4]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n22 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U6  ( .A1(
        CipherErrorVec2[5]), .A2(CipherErrorVec2[3]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n21 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U5  ( .A(Feedback[7]), 
        .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n20 ), .Z(Output[7])
         );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U4  ( .A1(
        CipherErrorVec2[3]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U3  ( .A1(
        CipherErrorVec2[5]), .A2(CipherErrorVec2[4]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n26 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U14  ( .A(Feedback[8]), 
        .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n27 ), .Z(Output[8])
         );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U13  ( .A1(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n26 ), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n27 ) );
  INV_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U12  ( .A(
        CipherErrorVec2[6]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U11  ( .A(Feedback[9]), 
        .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n24 ), .Z(Output[9])
         );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U10  ( .A1(
        CipherErrorVec2[8]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n23 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U9  ( .A1(
        CipherErrorVec2[7]), .A2(CipherErrorVec2[6]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n23 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U8  ( .A(Feedback[10]), 
        .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n22 ), .Z(Output[10])
         );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U7  ( .A1(
        CipherErrorVec2[7]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n22 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U6  ( .A1(
        CipherErrorVec2[8]), .A2(CipherErrorVec2[6]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n21 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U5  ( .A(Feedback[11]), 
        .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n20 ), .Z(Output[11])
         );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U4  ( .A1(
        CipherErrorVec2[6]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U3  ( .A1(
        CipherErrorVec2[8]), .A2(CipherErrorVec2[7]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n26 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U14  ( .A(
        Feedback[12]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n27 ), 
        .Z(Output[12]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U13  ( .A1(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n26 ), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n27 ) );
  INV_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U12  ( .A(
        CipherErrorVec2[9]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U11  ( .A(
        Feedback[13]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n24 ), 
        .Z(Output[13]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U10  ( .A1(
        CipherErrorVec2[11]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n23 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U9  ( .A1(
        CipherErrorVec2[10]), .A2(CipherErrorVec2[9]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n23 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U8  ( .A(Feedback[14]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n22 ), .Z(Output[14]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U7  ( .A1(
        CipherErrorVec2[10]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n22 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U6  ( .A1(
        CipherErrorVec2[11]), .A2(CipherErrorVec2[9]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n21 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U5  ( .A(Feedback[15]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n20 ), .Z(Output[15]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U4  ( .A1(
        CipherErrorVec2[9]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U3  ( .A1(
        CipherErrorVec2[11]), .A2(CipherErrorVec2[10]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n26 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U14  ( .A(
        Feedback[16]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n27 ), 
        .Z(Output[16]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U13  ( .A1(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n26 ), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n27 ) );
  INV_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U12  ( .A(
        CipherErrorVec2[12]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U11  ( .A(
        Feedback[17]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n24 ), 
        .Z(Output[17]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U10  ( .A1(
        CipherErrorVec2[14]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n23 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U9  ( .A1(
        CipherErrorVec2[13]), .A2(CipherErrorVec2[12]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n23 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U8  ( .A(Feedback[18]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n22 ), .Z(Output[18]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U7  ( .A1(
        CipherErrorVec2[13]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n22 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U6  ( .A1(
        CipherErrorVec2[14]), .A2(CipherErrorVec2[12]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n21 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U5  ( .A(Feedback[19]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n20 ), .Z(Output[19]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U4  ( .A1(
        CipherErrorVec2[12]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U3  ( .A1(
        CipherErrorVec2[14]), .A2(CipherErrorVec2[13]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n26 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U14  ( .A(
        Feedback[20]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n27 ), 
        .Z(Output[20]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U13  ( .A1(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n26 ), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n27 ) );
  INV_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U12  ( .A(
        CipherErrorVec2[15]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U11  ( .A(
        Feedback[21]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n24 ), 
        .Z(Output[21]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U10  ( .A1(
        CipherErrorVec2[17]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n23 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U9  ( .A1(
        CipherErrorVec2[16]), .A2(CipherErrorVec2[15]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n23 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U8  ( .A(Feedback[22]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n22 ), .Z(Output[22]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U7  ( .A1(
        CipherErrorVec2[16]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n22 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U6  ( .A1(
        CipherErrorVec2[17]), .A2(CipherErrorVec2[15]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n21 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U5  ( .A(Feedback[23]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n20 ), .Z(Output[23]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U4  ( .A1(
        CipherErrorVec2[15]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U3  ( .A1(
        CipherErrorVec2[17]), .A2(CipherErrorVec2[16]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n26 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U14  ( .A(
        Feedback[24]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n27 ), 
        .Z(Output[24]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U13  ( .A1(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n26 ), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n27 ) );
  INV_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U12  ( .A(
        CipherErrorVec2[18]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U11  ( .A(
        Feedback[25]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n24 ), 
        .Z(Output[25]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U10  ( .A1(
        CipherErrorVec2[20]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n23 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U9  ( .A1(
        CipherErrorVec2[19]), .A2(CipherErrorVec2[18]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n23 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U8  ( .A(Feedback[26]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n22 ), .Z(Output[26]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U7  ( .A1(
        CipherErrorVec2[19]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n22 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U6  ( .A1(
        CipherErrorVec2[20]), .A2(CipherErrorVec2[18]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n21 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U5  ( .A(Feedback[27]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n20 ), .Z(Output[27]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U4  ( .A1(
        CipherErrorVec2[18]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U3  ( .A1(
        CipherErrorVec2[20]), .A2(CipherErrorVec2[19]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n26 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U14  ( .A(
        Feedback[28]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n27 ), 
        .Z(Output[28]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U13  ( .A1(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n26 ), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n27 ) );
  INV_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U12  ( .A(
        CipherErrorVec2[21]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U11  ( .A(
        Feedback[29]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n24 ), 
        .Z(Output[29]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U10  ( .A1(
        CipherErrorVec2[23]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n23 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U9  ( .A1(
        CipherErrorVec2[22]), .A2(CipherErrorVec2[21]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n23 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U8  ( .A(Feedback[30]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n22 ), .Z(Output[30]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U7  ( .A1(
        CipherErrorVec2[22]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n22 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U6  ( .A1(
        CipherErrorVec2[23]), .A2(CipherErrorVec2[21]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n21 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U5  ( .A(Feedback[31]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n20 ), .Z(Output[31]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U4  ( .A1(
        CipherErrorVec2[21]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U3  ( .A1(
        CipherErrorVec2[23]), .A2(CipherErrorVec2[22]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n26 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U14  ( .A(
        Feedback[32]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n27 ), 
        .Z(Output[32]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U13  ( .A1(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n26 ), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n27 ) );
  INV_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U12  ( .A(
        CipherErrorVec2[24]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U11  ( .A(
        Feedback[33]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n24 ), 
        .Z(Output[33]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U10  ( .A1(
        CipherErrorVec2[26]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n23 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U9  ( .A1(
        CipherErrorVec2[25]), .A2(CipherErrorVec2[24]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n23 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U8  ( .A(Feedback[34]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n22 ), .Z(Output[34]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U7  ( .A1(
        CipherErrorVec2[25]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n22 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U6  ( .A1(
        CipherErrorVec2[26]), .A2(CipherErrorVec2[24]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n21 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U5  ( .A(Feedback[35]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n20 ), .Z(Output[35]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U4  ( .A1(
        CipherErrorVec2[24]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U3  ( .A1(
        CipherErrorVec2[26]), .A2(CipherErrorVec2[25]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n26 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U14  ( .A(
        Feedback[36]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n27 ), 
        .Z(Output[36]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U13  ( .A1(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n26 ), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n27 ) );
  INV_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U12  ( .A(
        CipherErrorVec2[27]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U11  ( .A(
        Feedback[37]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n24 ), 
        .Z(Output[37]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U10  ( .A1(
        CipherErrorVec2[29]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n23 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U9  ( .A1(
        CipherErrorVec2[28]), .A2(CipherErrorVec2[27]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n23 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U8  ( .A(Feedback[38]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n22 ), .Z(Output[38]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U7  ( .A1(
        CipherErrorVec2[28]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n22 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U6  ( .A1(
        CipherErrorVec2[29]), .A2(CipherErrorVec2[27]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n21 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U5  ( .A(Feedback[39]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n20 ), .Z(Output[39]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U4  ( .A1(
        CipherErrorVec2[27]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U3  ( .A1(
        CipherErrorVec2[29]), .A2(CipherErrorVec2[28]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n26 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U14  ( .A(
        Feedback[40]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n27 ), 
        .Z(Output[40]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U13  ( .A1(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n26 ), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n27 ) );
  INV_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U12  ( .A(
        CipherErrorVec2[30]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U11  ( .A(
        Feedback[41]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n24 ), 
        .Z(Output[41]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U10  ( .A1(
        CipherErrorVec2[32]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n23 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U9  ( .A1(
        CipherErrorVec2[31]), .A2(CipherErrorVec2[30]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n23 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U8  ( .A(Feedback[42]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n22 ), .Z(Output[42]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U7  ( .A1(
        CipherErrorVec2[31]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n22 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U6  ( .A1(
        CipherErrorVec2[32]), .A2(CipherErrorVec2[30]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n21 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U5  ( .A(Feedback[43]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n20 ), .Z(Output[43]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U4  ( .A1(
        CipherErrorVec2[30]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U3  ( .A1(
        CipherErrorVec2[32]), .A2(CipherErrorVec2[31]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n26 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U14  ( .A(
        Feedback[44]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n27 ), 
        .Z(Output[44]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U13  ( .A1(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n26 ), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n27 ) );
  INV_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U12  ( .A(
        CipherErrorVec2[33]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U11  ( .A(
        Feedback[45]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n24 ), 
        .Z(Output[45]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U10  ( .A1(
        CipherErrorVec2[35]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n23 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U9  ( .A1(
        CipherErrorVec2[34]), .A2(CipherErrorVec2[33]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n23 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U8  ( .A(Feedback[46]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n22 ), .Z(Output[46]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U7  ( .A1(
        CipherErrorVec2[34]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n22 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U6  ( .A1(
        CipherErrorVec2[35]), .A2(CipherErrorVec2[33]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n21 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U5  ( .A(Feedback[47]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n20 ), .Z(Output[47]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U4  ( .A1(
        CipherErrorVec2[33]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U3  ( .A1(
        CipherErrorVec2[35]), .A2(CipherErrorVec2[34]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n26 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U14  ( .A(
        Feedback[48]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n27 ), 
        .Z(Output[48]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U13  ( .A1(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n26 ), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n27 ) );
  INV_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U12  ( .A(
        CipherErrorVec2[36]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U11  ( .A(
        Feedback[49]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n24 ), 
        .Z(Output[49]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U10  ( .A1(
        CipherErrorVec2[38]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n23 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U9  ( .A1(
        CipherErrorVec2[37]), .A2(CipherErrorVec2[36]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n23 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U8  ( .A(Feedback[50]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n22 ), .Z(Output[50]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U7  ( .A1(
        CipherErrorVec2[37]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n22 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U6  ( .A1(
        CipherErrorVec2[38]), .A2(CipherErrorVec2[36]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n21 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U5  ( .A(Feedback[51]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n20 ), .Z(Output[51]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U4  ( .A1(
        CipherErrorVec2[36]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U3  ( .A1(
        CipherErrorVec2[38]), .A2(CipherErrorVec2[37]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n26 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U14  ( .A(
        Feedback[52]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n27 ), 
        .Z(Output[52]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U13  ( .A1(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n26 ), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n27 ) );
  INV_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U12  ( .A(
        CipherErrorVec2[39]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U11  ( .A(
        Feedback[53]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n24 ), 
        .Z(Output[53]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U10  ( .A1(
        CipherErrorVec2[41]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n23 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U9  ( .A1(
        CipherErrorVec2[40]), .A2(CipherErrorVec2[39]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n23 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U8  ( .A(Feedback[54]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n22 ), .Z(Output[54]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U7  ( .A1(
        CipherErrorVec2[40]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n22 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U6  ( .A1(
        CipherErrorVec2[41]), .A2(CipherErrorVec2[39]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n21 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U5  ( .A(Feedback[55]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n20 ), .Z(Output[55]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U4  ( .A1(
        CipherErrorVec2[39]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U3  ( .A1(
        CipherErrorVec2[41]), .A2(CipherErrorVec2[40]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n26 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U14  ( .A(
        Feedback[56]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n27 ), 
        .Z(Output[56]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U13  ( .A1(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n26 ), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n27 ) );
  INV_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U12  ( .A(
        CipherErrorVec2[42]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U11  ( .A(
        Feedback[57]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n24 ), 
        .Z(Output[57]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U10  ( .A1(
        CipherErrorVec2[44]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n23 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U9  ( .A1(
        CipherErrorVec2[43]), .A2(CipherErrorVec2[42]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n23 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U8  ( .A(Feedback[58]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n22 ), .Z(Output[58]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U7  ( .A1(
        CipherErrorVec2[43]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n22 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U6  ( .A1(
        CipherErrorVec2[44]), .A2(CipherErrorVec2[42]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n21 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U5  ( .A(Feedback[59]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n20 ), .Z(Output[59]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U4  ( .A1(
        CipherErrorVec2[42]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U3  ( .A1(
        CipherErrorVec2[44]), .A2(CipherErrorVec2[43]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n26 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U14  ( .A(
        Feedback[60]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n27 ), 
        .Z(Output[60]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U13  ( .A1(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n26 ), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n25 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n27 ) );
  INV_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U12  ( .A(
        CipherErrorVec2[45]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n25 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U11  ( .A(
        Feedback[61]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n24 ), 
        .Z(Output[61]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U10  ( .A1(
        CipherErrorVec2[47]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n23 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n24 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U9  ( .A1(
        CipherErrorVec2[46]), .A2(CipherErrorVec2[45]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n23 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U8  ( .A(Feedback[62]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n22 ), .Z(Output[62]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U7  ( .A1(
        CipherErrorVec2[46]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n21 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n22 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U6  ( .A1(
        CipherErrorVec2[47]), .A2(CipherErrorVec2[45]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n21 ) );
  XOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U5  ( .A(Feedback[63]), .B(\SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n20 ), .Z(Output[63]) );
  NOR2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U4  ( .A1(
        CipherErrorVec2[45]), .A2(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n26 ), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n20 ) );
  NAND2_X1 \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U3  ( .A1(
        CipherErrorVec2[47]), .A2(CipherErrorVec2[46]), .ZN(
        \SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n26 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_0_LFInst_0_n2 ), .B(Key[1]), .ZN(Red_K0[0]) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_0_U3  ( .A(Key[2]), .B(Key[0]), .ZN(
        \Red_K0Inst_LFInst_0_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_0_LFInst_1_n2 ), .B(Key[1]), .ZN(Red_K0[1]) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_1_U3  ( .A(Key[3]), .B(Key[0]), .ZN(
        \Red_K0Inst_LFInst_0_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_0_LFInst_2_n2 ), .B(Key[2]), .ZN(Red_K0[2]) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_2_U3  ( .A(Key[3]), .B(Key[0]), .ZN(
        \Red_K0Inst_LFInst_0_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_1_LFInst_0_n2 ), .B(Key[5]), .ZN(Red_K0[3]) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_0_U3  ( .A(Key[6]), .B(Key[4]), .ZN(
        \Red_K0Inst_LFInst_1_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_1_LFInst_1_n2 ), .B(Key[5]), .ZN(Red_K0[4]) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_1_U3  ( .A(Key[7]), .B(Key[4]), .ZN(
        \Red_K0Inst_LFInst_1_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_1_LFInst_2_n2 ), .B(Key[6]), .ZN(Red_K0[5]) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_2_U3  ( .A(Key[7]), .B(Key[4]), .ZN(
        \Red_K0Inst_LFInst_1_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_2_LFInst_0_n2 ), .B(Key[9]), .ZN(Red_K0[6]) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_0_U3  ( .A(Key[10]), .B(Key[8]), .ZN(
        \Red_K0Inst_LFInst_2_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_2_LFInst_1_n2 ), .B(Key[9]), .ZN(Red_K0[7]) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_1_U3  ( .A(Key[11]), .B(Key[8]), .ZN(
        \Red_K0Inst_LFInst_2_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_2_LFInst_2_n2 ), .B(Key[10]), .ZN(Red_K0[8]) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_2_U3  ( .A(Key[11]), .B(Key[8]), .ZN(
        \Red_K0Inst_LFInst_2_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_3_LFInst_0_n2 ), .B(Key[13]), .ZN(Red_K0[9]) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_0_U3  ( .A(Key[14]), .B(Key[12]), .ZN(
        \Red_K0Inst_LFInst_3_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_3_LFInst_1_n2 ), .B(Key[13]), .ZN(Red_K0[10]) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_1_U3  ( .A(Key[15]), .B(Key[12]), .ZN(
        \Red_K0Inst_LFInst_3_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_3_LFInst_2_n2 ), .B(Key[14]), .ZN(Red_K0[11]) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_2_U3  ( .A(Key[15]), .B(Key[12]), .ZN(
        \Red_K0Inst_LFInst_3_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_4_LFInst_0_n2 ), .B(Key[17]), .ZN(Red_K0[12]) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_0_U3  ( .A(Key[18]), .B(Key[16]), .ZN(
        \Red_K0Inst_LFInst_4_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_4_LFInst_1_n2 ), .B(Key[17]), .ZN(Red_K0[13]) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_1_U3  ( .A(Key[19]), .B(Key[16]), .ZN(
        \Red_K0Inst_LFInst_4_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_4_LFInst_2_n2 ), .B(Key[18]), .ZN(Red_K0[14]) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_2_U3  ( .A(Key[19]), .B(Key[16]), .ZN(
        \Red_K0Inst_LFInst_4_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_5_LFInst_0_n2 ), .B(Key[21]), .ZN(Red_K0[15]) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_0_U3  ( .A(Key[22]), .B(Key[20]), .ZN(
        \Red_K0Inst_LFInst_5_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_5_LFInst_1_n2 ), .B(Key[21]), .ZN(Red_K0[16]) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_1_U3  ( .A(Key[23]), .B(Key[20]), .ZN(
        \Red_K0Inst_LFInst_5_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_5_LFInst_2_n2 ), .B(Key[22]), .ZN(Red_K0[17]) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_2_U3  ( .A(Key[23]), .B(Key[20]), .ZN(
        \Red_K0Inst_LFInst_5_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_6_LFInst_0_n2 ), .B(Key[25]), .ZN(Red_K0[18]) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_0_U3  ( .A(Key[26]), .B(Key[24]), .ZN(
        \Red_K0Inst_LFInst_6_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_6_LFInst_1_n2 ), .B(Key[25]), .ZN(Red_K0[19]) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_1_U3  ( .A(Key[27]), .B(Key[24]), .ZN(
        \Red_K0Inst_LFInst_6_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_6_LFInst_2_n2 ), .B(Key[26]), .ZN(Red_K0[20]) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_2_U3  ( .A(Key[27]), .B(Key[24]), .ZN(
        \Red_K0Inst_LFInst_6_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_7_LFInst_0_n2 ), .B(Key[29]), .ZN(Red_K0[21]) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_0_U3  ( .A(Key[30]), .B(Key[28]), .ZN(
        \Red_K0Inst_LFInst_7_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_7_LFInst_1_n2 ), .B(Key[29]), .ZN(Red_K0[22]) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_1_U3  ( .A(Key[31]), .B(Key[28]), .ZN(
        \Red_K0Inst_LFInst_7_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_7_LFInst_2_n2 ), .B(Key[30]), .ZN(Red_K0[23]) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_2_U3  ( .A(Key[31]), .B(Key[28]), .ZN(
        \Red_K0Inst_LFInst_7_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_8_LFInst_0_n2 ), .B(Key[33]), .ZN(Red_K0[24]) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_0_U3  ( .A(Key[34]), .B(Key[32]), .ZN(
        \Red_K0Inst_LFInst_8_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_8_LFInst_1_n2 ), .B(Key[33]), .ZN(Red_K0[25]) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_1_U3  ( .A(Key[35]), .B(Key[32]), .ZN(
        \Red_K0Inst_LFInst_8_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_8_LFInst_2_n2 ), .B(Key[34]), .ZN(Red_K0[26]) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_2_U3  ( .A(Key[35]), .B(Key[32]), .ZN(
        \Red_K0Inst_LFInst_8_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_9_LFInst_0_n2 ), .B(Key[37]), .ZN(Red_K0[27]) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_0_U3  ( .A(Key[38]), .B(Key[36]), .ZN(
        \Red_K0Inst_LFInst_9_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_9_LFInst_1_n2 ), .B(Key[37]), .ZN(Red_K0[28]) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_1_U3  ( .A(Key[39]), .B(Key[36]), .ZN(
        \Red_K0Inst_LFInst_9_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_9_LFInst_2_n2 ), .B(Key[38]), .ZN(Red_K0[29]) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_2_U3  ( .A(Key[39]), .B(Key[36]), .ZN(
        \Red_K0Inst_LFInst_9_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_10_LFInst_0_n2 ), .B(Key[41]), .ZN(Red_K0[30]) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_0_U3  ( .A(Key[42]), .B(Key[40]), .ZN(
        \Red_K0Inst_LFInst_10_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_10_LFInst_1_n2 ), .B(Key[41]), .ZN(Red_K0[31]) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_1_U3  ( .A(Key[43]), .B(Key[40]), .ZN(
        \Red_K0Inst_LFInst_10_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_10_LFInst_2_n2 ), .B(Key[42]), .ZN(Red_K0[32]) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_2_U3  ( .A(Key[43]), .B(Key[40]), .ZN(
        \Red_K0Inst_LFInst_10_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_11_LFInst_0_n2 ), .B(Key[45]), .ZN(Red_K0[33]) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_0_U3  ( .A(Key[46]), .B(Key[44]), .ZN(
        \Red_K0Inst_LFInst_11_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_11_LFInst_1_n2 ), .B(Key[45]), .ZN(Red_K0[34]) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_1_U3  ( .A(Key[47]), .B(Key[44]), .ZN(
        \Red_K0Inst_LFInst_11_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_11_LFInst_2_n2 ), .B(Key[46]), .ZN(Red_K0[35]) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_2_U3  ( .A(Key[47]), .B(Key[44]), .ZN(
        \Red_K0Inst_LFInst_11_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_12_LFInst_0_n2 ), .B(Key[49]), .ZN(Red_K0[36]) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_0_U3  ( .A(Key[50]), .B(Key[48]), .ZN(
        \Red_K0Inst_LFInst_12_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_12_LFInst_1_n2 ), .B(Key[49]), .ZN(Red_K0[37]) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_1_U3  ( .A(Key[51]), .B(Key[48]), .ZN(
        \Red_K0Inst_LFInst_12_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_12_LFInst_2_n2 ), .B(Key[50]), .ZN(Red_K0[38]) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_2_U3  ( .A(Key[51]), .B(Key[48]), .ZN(
        \Red_K0Inst_LFInst_12_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_13_LFInst_0_n2 ), .B(Key[53]), .ZN(Red_K0[39]) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_0_U3  ( .A(Key[54]), .B(Key[52]), .ZN(
        \Red_K0Inst_LFInst_13_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_13_LFInst_1_n2 ), .B(Key[53]), .ZN(Red_K0[40]) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_1_U3  ( .A(Key[55]), .B(Key[52]), .ZN(
        \Red_K0Inst_LFInst_13_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_13_LFInst_2_n2 ), .B(Key[54]), .ZN(Red_K0[41]) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_2_U3  ( .A(Key[55]), .B(Key[52]), .ZN(
        \Red_K0Inst_LFInst_13_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_14_LFInst_0_n2 ), .B(Key[57]), .ZN(Red_K0[42]) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_0_U3  ( .A(Key[58]), .B(Key[56]), .ZN(
        \Red_K0Inst_LFInst_14_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_14_LFInst_1_n2 ), .B(Key[57]), .ZN(Red_K0[43]) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_1_U3  ( .A(Key[59]), .B(Key[56]), .ZN(
        \Red_K0Inst_LFInst_14_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_14_LFInst_2_n2 ), .B(Key[58]), .ZN(Red_K0[44]) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_2_U3  ( .A(Key[59]), .B(Key[56]), .ZN(
        \Red_K0Inst_LFInst_14_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_15_LFInst_0_n2 ), .B(Key[61]), .ZN(Red_K0[45]) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_0_U3  ( .A(Key[62]), .B(Key[60]), .ZN(
        \Red_K0Inst_LFInst_15_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_15_LFInst_1_n2 ), .B(Key[61]), .ZN(Red_K0[46]) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_1_U3  ( .A(Key[63]), .B(Key[60]), .ZN(
        \Red_K0Inst_LFInst_15_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_15_LFInst_2_n2 ), .B(Key[62]), .ZN(Red_K0[47]) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_2_U3  ( .A(Key[63]), .B(Key[60]), .ZN(
        \Red_K0Inst_LFInst_15_LFInst_2_n2 ) );
endmodule

