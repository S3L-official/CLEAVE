module LED64Enc ( clk, rst, Plaintext, Key, Ciphertext, ErrorFlag );
  input [63:0] Plaintext;
  input [63:0] Key;
  output [63:0] Ciphertext;
  (* FIRMER="clock" *)input clk, rst;
  output ErrorFlag;
  wire   n5, \SubCellInst_LFInst_0_LFInst_0_n9 ,
         \SubCellInst_LFInst_0_LFInst_0_n8 ,
         \SubCellInst_LFInst_0_LFInst_0_n7 ,
         \SubCellInst_LFInst_0_LFInst_0_n10 ,
         \SubCellInst_LFInst_0_LFInst_1_n18 ,
         \SubCellInst_LFInst_0_LFInst_1_n17 ,
         \SubCellInst_LFInst_0_LFInst_1_n16 ,
         \SubCellInst_LFInst_0_LFInst_1_n15 ,
         \SubCellInst_LFInst_0_LFInst_1_n14 ,
         \SubCellInst_LFInst_0_LFInst_1_n13 ,
         \SubCellInst_LFInst_0_LFInst_1_n12 ,
         \SubCellInst_LFInst_0_LFInst_1_n11 ,
         \SubCellInst_LFInst_0_LFInst_1_n10 ,
         \SubCellInst_LFInst_0_LFInst_2_n22 ,
         \SubCellInst_LFInst_0_LFInst_2_n21 ,
         \SubCellInst_LFInst_0_LFInst_2_n20 ,
         \SubCellInst_LFInst_0_LFInst_2_n19 ,
         \SubCellInst_LFInst_0_LFInst_2_n18 ,
         \SubCellInst_LFInst_0_LFInst_2_n17 ,
         \SubCellInst_LFInst_0_LFInst_2_n16 ,
         \SubCellInst_LFInst_0_LFInst_2_n15 ,
         \SubCellInst_LFInst_0_LFInst_3_n16 ,
         \SubCellInst_LFInst_0_LFInst_3_n15 ,
         \SubCellInst_LFInst_0_LFInst_3_n14 ,
         \SubCellInst_LFInst_0_LFInst_3_n13 ,
         \SubCellInst_LFInst_0_LFInst_3_n12 ,
         \SubCellInst_LFInst_0_LFInst_3_n11 ,
         \SubCellInst_LFInst_1_LFInst_0_n10 ,
         \SubCellInst_LFInst_1_LFInst_0_n9 ,
         \SubCellInst_LFInst_1_LFInst_0_n8 ,
         \SubCellInst_LFInst_1_LFInst_0_n7 ,
         \SubCellInst_LFInst_1_LFInst_1_n18 ,
         \SubCellInst_LFInst_1_LFInst_1_n17 ,
         \SubCellInst_LFInst_1_LFInst_1_n16 ,
         \SubCellInst_LFInst_1_LFInst_1_n15 ,
         \SubCellInst_LFInst_1_LFInst_1_n14 ,
         \SubCellInst_LFInst_1_LFInst_1_n13 ,
         \SubCellInst_LFInst_1_LFInst_1_n12 ,
         \SubCellInst_LFInst_1_LFInst_1_n11 ,
         \SubCellInst_LFInst_1_LFInst_1_n10 ,
         \SubCellInst_LFInst_1_LFInst_2_n22 ,
         \SubCellInst_LFInst_1_LFInst_2_n21 ,
         \SubCellInst_LFInst_1_LFInst_2_n20 ,
         \SubCellInst_LFInst_1_LFInst_2_n19 ,
         \SubCellInst_LFInst_1_LFInst_2_n18 ,
         \SubCellInst_LFInst_1_LFInst_2_n17 ,
         \SubCellInst_LFInst_1_LFInst_2_n16 ,
         \SubCellInst_LFInst_1_LFInst_2_n15 ,
         \SubCellInst_LFInst_1_LFInst_3_n16 ,
         \SubCellInst_LFInst_1_LFInst_3_n15 ,
         \SubCellInst_LFInst_1_LFInst_3_n14 ,
         \SubCellInst_LFInst_1_LFInst_3_n13 ,
         \SubCellInst_LFInst_1_LFInst_3_n12 ,
         \SubCellInst_LFInst_1_LFInst_3_n11 ,
         \SubCellInst_LFInst_2_LFInst_0_n10 ,
         \SubCellInst_LFInst_2_LFInst_0_n9 ,
         \SubCellInst_LFInst_2_LFInst_0_n8 ,
         \SubCellInst_LFInst_2_LFInst_0_n7 ,
         \SubCellInst_LFInst_2_LFInst_1_n18 ,
         \SubCellInst_LFInst_2_LFInst_1_n17 ,
         \SubCellInst_LFInst_2_LFInst_1_n16 ,
         \SubCellInst_LFInst_2_LFInst_1_n15 ,
         \SubCellInst_LFInst_2_LFInst_1_n14 ,
         \SubCellInst_LFInst_2_LFInst_1_n13 ,
         \SubCellInst_LFInst_2_LFInst_1_n12 ,
         \SubCellInst_LFInst_2_LFInst_1_n11 ,
         \SubCellInst_LFInst_2_LFInst_1_n10 ,
         \SubCellInst_LFInst_2_LFInst_2_n22 ,
         \SubCellInst_LFInst_2_LFInst_2_n21 ,
         \SubCellInst_LFInst_2_LFInst_2_n20 ,
         \SubCellInst_LFInst_2_LFInst_2_n19 ,
         \SubCellInst_LFInst_2_LFInst_2_n18 ,
         \SubCellInst_LFInst_2_LFInst_2_n17 ,
         \SubCellInst_LFInst_2_LFInst_2_n16 ,
         \SubCellInst_LFInst_2_LFInst_2_n15 ,
         \SubCellInst_LFInst_2_LFInst_3_n16 ,
         \SubCellInst_LFInst_2_LFInst_3_n15 ,
         \SubCellInst_LFInst_2_LFInst_3_n14 ,
         \SubCellInst_LFInst_2_LFInst_3_n13 ,
         \SubCellInst_LFInst_2_LFInst_3_n12 ,
         \SubCellInst_LFInst_2_LFInst_3_n11 ,
         \SubCellInst_LFInst_3_LFInst_0_n10 ,
         \SubCellInst_LFInst_3_LFInst_0_n9 ,
         \SubCellInst_LFInst_3_LFInst_0_n8 ,
         \SubCellInst_LFInst_3_LFInst_0_n7 ,
         \SubCellInst_LFInst_3_LFInst_1_n18 ,
         \SubCellInst_LFInst_3_LFInst_1_n17 ,
         \SubCellInst_LFInst_3_LFInst_1_n16 ,
         \SubCellInst_LFInst_3_LFInst_1_n15 ,
         \SubCellInst_LFInst_3_LFInst_1_n14 ,
         \SubCellInst_LFInst_3_LFInst_1_n13 ,
         \SubCellInst_LFInst_3_LFInst_1_n12 ,
         \SubCellInst_LFInst_3_LFInst_1_n11 ,
         \SubCellInst_LFInst_3_LFInst_1_n10 ,
         \SubCellInst_LFInst_3_LFInst_2_n22 ,
         \SubCellInst_LFInst_3_LFInst_2_n21 ,
         \SubCellInst_LFInst_3_LFInst_2_n20 ,
         \SubCellInst_LFInst_3_LFInst_2_n19 ,
         \SubCellInst_LFInst_3_LFInst_2_n18 ,
         \SubCellInst_LFInst_3_LFInst_2_n17 ,
         \SubCellInst_LFInst_3_LFInst_2_n16 ,
         \SubCellInst_LFInst_3_LFInst_2_n15 ,
         \SubCellInst_LFInst_3_LFInst_3_n16 ,
         \SubCellInst_LFInst_3_LFInst_3_n15 ,
         \SubCellInst_LFInst_3_LFInst_3_n14 ,
         \SubCellInst_LFInst_3_LFInst_3_n13 ,
         \SubCellInst_LFInst_3_LFInst_3_n12 ,
         \SubCellInst_LFInst_3_LFInst_3_n11 ,
         \SubCellInst_LFInst_4_LFInst_0_n9 ,
         \SubCellInst_LFInst_4_LFInst_0_n8 ,
         \SubCellInst_LFInst_4_LFInst_0_n7 ,
         \SubCellInst_LFInst_4_LFInst_0_n10 ,
         \SubCellInst_LFInst_4_LFInst_1_n18 ,
         \SubCellInst_LFInst_4_LFInst_1_n17 ,
         \SubCellInst_LFInst_4_LFInst_1_n16 ,
         \SubCellInst_LFInst_4_LFInst_1_n15 ,
         \SubCellInst_LFInst_4_LFInst_1_n14 ,
         \SubCellInst_LFInst_4_LFInst_1_n13 ,
         \SubCellInst_LFInst_4_LFInst_1_n12 ,
         \SubCellInst_LFInst_4_LFInst_1_n11 ,
         \SubCellInst_LFInst_4_LFInst_1_n10 ,
         \SubCellInst_LFInst_4_LFInst_2_n22 ,
         \SubCellInst_LFInst_4_LFInst_2_n21 ,
         \SubCellInst_LFInst_4_LFInst_2_n20 ,
         \SubCellInst_LFInst_4_LFInst_2_n19 ,
         \SubCellInst_LFInst_4_LFInst_2_n18 ,
         \SubCellInst_LFInst_4_LFInst_2_n17 ,
         \SubCellInst_LFInst_4_LFInst_2_n16 ,
         \SubCellInst_LFInst_4_LFInst_2_n15 ,
         \SubCellInst_LFInst_4_LFInst_3_n16 ,
         \SubCellInst_LFInst_4_LFInst_3_n15 ,
         \SubCellInst_LFInst_4_LFInst_3_n14 ,
         \SubCellInst_LFInst_4_LFInst_3_n13 ,
         \SubCellInst_LFInst_4_LFInst_3_n12 ,
         \SubCellInst_LFInst_4_LFInst_3_n11 ,
         \SubCellInst_LFInst_5_LFInst_0_n10 ,
         \SubCellInst_LFInst_5_LFInst_0_n9 ,
         \SubCellInst_LFInst_5_LFInst_0_n8 ,
         \SubCellInst_LFInst_5_LFInst_0_n7 ,
         \SubCellInst_LFInst_5_LFInst_1_n18 ,
         \SubCellInst_LFInst_5_LFInst_1_n17 ,
         \SubCellInst_LFInst_5_LFInst_1_n16 ,
         \SubCellInst_LFInst_5_LFInst_1_n15 ,
         \SubCellInst_LFInst_5_LFInst_1_n14 ,
         \SubCellInst_LFInst_5_LFInst_1_n13 ,
         \SubCellInst_LFInst_5_LFInst_1_n12 ,
         \SubCellInst_LFInst_5_LFInst_1_n11 ,
         \SubCellInst_LFInst_5_LFInst_1_n10 ,
         \SubCellInst_LFInst_5_LFInst_2_n22 ,
         \SubCellInst_LFInst_5_LFInst_2_n21 ,
         \SubCellInst_LFInst_5_LFInst_2_n20 ,
         \SubCellInst_LFInst_5_LFInst_2_n19 ,
         \SubCellInst_LFInst_5_LFInst_2_n18 ,
         \SubCellInst_LFInst_5_LFInst_2_n17 ,
         \SubCellInst_LFInst_5_LFInst_2_n16 ,
         \SubCellInst_LFInst_5_LFInst_2_n15 ,
         \SubCellInst_LFInst_5_LFInst_3_n16 ,
         \SubCellInst_LFInst_5_LFInst_3_n15 ,
         \SubCellInst_LFInst_5_LFInst_3_n14 ,
         \SubCellInst_LFInst_5_LFInst_3_n13 ,
         \SubCellInst_LFInst_5_LFInst_3_n12 ,
         \SubCellInst_LFInst_5_LFInst_3_n11 ,
         \SubCellInst_LFInst_6_LFInst_0_n10 ,
         \SubCellInst_LFInst_6_LFInst_0_n9 ,
         \SubCellInst_LFInst_6_LFInst_0_n8 ,
         \SubCellInst_LFInst_6_LFInst_0_n7 ,
         \SubCellInst_LFInst_6_LFInst_1_n18 ,
         \SubCellInst_LFInst_6_LFInst_1_n17 ,
         \SubCellInst_LFInst_6_LFInst_1_n16 ,
         \SubCellInst_LFInst_6_LFInst_1_n15 ,
         \SubCellInst_LFInst_6_LFInst_1_n14 ,
         \SubCellInst_LFInst_6_LFInst_1_n13 ,
         \SubCellInst_LFInst_6_LFInst_1_n12 ,
         \SubCellInst_LFInst_6_LFInst_1_n11 ,
         \SubCellInst_LFInst_6_LFInst_1_n10 ,
         \SubCellInst_LFInst_6_LFInst_2_n22 ,
         \SubCellInst_LFInst_6_LFInst_2_n21 ,
         \SubCellInst_LFInst_6_LFInst_2_n20 ,
         \SubCellInst_LFInst_6_LFInst_2_n19 ,
         \SubCellInst_LFInst_6_LFInst_2_n18 ,
         \SubCellInst_LFInst_6_LFInst_2_n17 ,
         \SubCellInst_LFInst_6_LFInst_2_n16 ,
         \SubCellInst_LFInst_6_LFInst_2_n15 ,
         \SubCellInst_LFInst_6_LFInst_3_n16 ,
         \SubCellInst_LFInst_6_LFInst_3_n15 ,
         \SubCellInst_LFInst_6_LFInst_3_n14 ,
         \SubCellInst_LFInst_6_LFInst_3_n13 ,
         \SubCellInst_LFInst_6_LFInst_3_n12 ,
         \SubCellInst_LFInst_6_LFInst_3_n11 ,
         \SubCellInst_LFInst_7_LFInst_0_n10 ,
         \SubCellInst_LFInst_7_LFInst_0_n9 ,
         \SubCellInst_LFInst_7_LFInst_0_n8 ,
         \SubCellInst_LFInst_7_LFInst_0_n7 ,
         \SubCellInst_LFInst_7_LFInst_1_n18 ,
         \SubCellInst_LFInst_7_LFInst_1_n17 ,
         \SubCellInst_LFInst_7_LFInst_1_n16 ,
         \SubCellInst_LFInst_7_LFInst_1_n15 ,
         \SubCellInst_LFInst_7_LFInst_1_n14 ,
         \SubCellInst_LFInst_7_LFInst_1_n13 ,
         \SubCellInst_LFInst_7_LFInst_1_n12 ,
         \SubCellInst_LFInst_7_LFInst_1_n11 ,
         \SubCellInst_LFInst_7_LFInst_1_n10 ,
         \SubCellInst_LFInst_7_LFInst_2_n22 ,
         \SubCellInst_LFInst_7_LFInst_2_n21 ,
         \SubCellInst_LFInst_7_LFInst_2_n20 ,
         \SubCellInst_LFInst_7_LFInst_2_n19 ,
         \SubCellInst_LFInst_7_LFInst_2_n18 ,
         \SubCellInst_LFInst_7_LFInst_2_n17 ,
         \SubCellInst_LFInst_7_LFInst_2_n16 ,
         \SubCellInst_LFInst_7_LFInst_2_n15 ,
         \SubCellInst_LFInst_7_LFInst_3_n16 ,
         \SubCellInst_LFInst_7_LFInst_3_n15 ,
         \SubCellInst_LFInst_7_LFInst_3_n14 ,
         \SubCellInst_LFInst_7_LFInst_3_n13 ,
         \SubCellInst_LFInst_7_LFInst_3_n12 ,
         \SubCellInst_LFInst_7_LFInst_3_n11 ,
         \SubCellInst_LFInst_8_LFInst_0_n10 ,
         \SubCellInst_LFInst_8_LFInst_0_n9 ,
         \SubCellInst_LFInst_8_LFInst_0_n8 ,
         \SubCellInst_LFInst_8_LFInst_0_n7 ,
         \SubCellInst_LFInst_8_LFInst_1_n18 ,
         \SubCellInst_LFInst_8_LFInst_1_n17 ,
         \SubCellInst_LFInst_8_LFInst_1_n16 ,
         \SubCellInst_LFInst_8_LFInst_1_n15 ,
         \SubCellInst_LFInst_8_LFInst_1_n14 ,
         \SubCellInst_LFInst_8_LFInst_1_n13 ,
         \SubCellInst_LFInst_8_LFInst_1_n12 ,
         \SubCellInst_LFInst_8_LFInst_1_n11 ,
         \SubCellInst_LFInst_8_LFInst_1_n10 ,
         \SubCellInst_LFInst_8_LFInst_2_n22 ,
         \SubCellInst_LFInst_8_LFInst_2_n21 ,
         \SubCellInst_LFInst_8_LFInst_2_n20 ,
         \SubCellInst_LFInst_8_LFInst_2_n19 ,
         \SubCellInst_LFInst_8_LFInst_2_n18 ,
         \SubCellInst_LFInst_8_LFInst_2_n17 ,
         \SubCellInst_LFInst_8_LFInst_2_n16 ,
         \SubCellInst_LFInst_8_LFInst_2_n15 ,
         \SubCellInst_LFInst_8_LFInst_3_n16 ,
         \SubCellInst_LFInst_8_LFInst_3_n15 ,
         \SubCellInst_LFInst_8_LFInst_3_n14 ,
         \SubCellInst_LFInst_8_LFInst_3_n13 ,
         \SubCellInst_LFInst_8_LFInst_3_n12 ,
         \SubCellInst_LFInst_8_LFInst_3_n11 ,
         \SubCellInst_LFInst_9_LFInst_0_n10 ,
         \SubCellInst_LFInst_9_LFInst_0_n9 ,
         \SubCellInst_LFInst_9_LFInst_0_n8 ,
         \SubCellInst_LFInst_9_LFInst_0_n7 ,
         \SubCellInst_LFInst_9_LFInst_1_n18 ,
         \SubCellInst_LFInst_9_LFInst_1_n17 ,
         \SubCellInst_LFInst_9_LFInst_1_n16 ,
         \SubCellInst_LFInst_9_LFInst_1_n15 ,
         \SubCellInst_LFInst_9_LFInst_1_n14 ,
         \SubCellInst_LFInst_9_LFInst_1_n13 ,
         \SubCellInst_LFInst_9_LFInst_1_n12 ,
         \SubCellInst_LFInst_9_LFInst_1_n11 ,
         \SubCellInst_LFInst_9_LFInst_1_n10 ,
         \SubCellInst_LFInst_9_LFInst_2_n22 ,
         \SubCellInst_LFInst_9_LFInst_2_n21 ,
         \SubCellInst_LFInst_9_LFInst_2_n20 ,
         \SubCellInst_LFInst_9_LFInst_2_n19 ,
         \SubCellInst_LFInst_9_LFInst_2_n18 ,
         \SubCellInst_LFInst_9_LFInst_2_n17 ,
         \SubCellInst_LFInst_9_LFInst_2_n16 ,
         \SubCellInst_LFInst_9_LFInst_2_n15 ,
         \SubCellInst_LFInst_9_LFInst_3_n16 ,
         \SubCellInst_LFInst_9_LFInst_3_n15 ,
         \SubCellInst_LFInst_9_LFInst_3_n14 ,
         \SubCellInst_LFInst_9_LFInst_3_n13 ,
         \SubCellInst_LFInst_9_LFInst_3_n12 ,
         \SubCellInst_LFInst_9_LFInst_3_n11 ,
         \SubCellInst_LFInst_10_LFInst_0_n10 ,
         \SubCellInst_LFInst_10_LFInst_0_n9 ,
         \SubCellInst_LFInst_10_LFInst_0_n8 ,
         \SubCellInst_LFInst_10_LFInst_0_n7 ,
         \SubCellInst_LFInst_10_LFInst_1_n18 ,
         \SubCellInst_LFInst_10_LFInst_1_n17 ,
         \SubCellInst_LFInst_10_LFInst_1_n16 ,
         \SubCellInst_LFInst_10_LFInst_1_n15 ,
         \SubCellInst_LFInst_10_LFInst_1_n14 ,
         \SubCellInst_LFInst_10_LFInst_1_n13 ,
         \SubCellInst_LFInst_10_LFInst_1_n12 ,
         \SubCellInst_LFInst_10_LFInst_1_n11 ,
         \SubCellInst_LFInst_10_LFInst_1_n10 ,
         \SubCellInst_LFInst_10_LFInst_2_n22 ,
         \SubCellInst_LFInst_10_LFInst_2_n21 ,
         \SubCellInst_LFInst_10_LFInst_2_n20 ,
         \SubCellInst_LFInst_10_LFInst_2_n19 ,
         \SubCellInst_LFInst_10_LFInst_2_n18 ,
         \SubCellInst_LFInst_10_LFInst_2_n17 ,
         \SubCellInst_LFInst_10_LFInst_2_n16 ,
         \SubCellInst_LFInst_10_LFInst_2_n15 ,
         \SubCellInst_LFInst_10_LFInst_3_n16 ,
         \SubCellInst_LFInst_10_LFInst_3_n15 ,
         \SubCellInst_LFInst_10_LFInst_3_n14 ,
         \SubCellInst_LFInst_10_LFInst_3_n13 ,
         \SubCellInst_LFInst_10_LFInst_3_n12 ,
         \SubCellInst_LFInst_10_LFInst_3_n11 ,
         \SubCellInst_LFInst_11_LFInst_0_n10 ,
         \SubCellInst_LFInst_11_LFInst_0_n9 ,
         \SubCellInst_LFInst_11_LFInst_0_n8 ,
         \SubCellInst_LFInst_11_LFInst_0_n7 ,
         \SubCellInst_LFInst_11_LFInst_1_n18 ,
         \SubCellInst_LFInst_11_LFInst_1_n17 ,
         \SubCellInst_LFInst_11_LFInst_1_n16 ,
         \SubCellInst_LFInst_11_LFInst_1_n15 ,
         \SubCellInst_LFInst_11_LFInst_1_n14 ,
         \SubCellInst_LFInst_11_LFInst_1_n13 ,
         \SubCellInst_LFInst_11_LFInst_1_n12 ,
         \SubCellInst_LFInst_11_LFInst_1_n11 ,
         \SubCellInst_LFInst_11_LFInst_1_n10 ,
         \SubCellInst_LFInst_11_LFInst_2_n22 ,
         \SubCellInst_LFInst_11_LFInst_2_n21 ,
         \SubCellInst_LFInst_11_LFInst_2_n20 ,
         \SubCellInst_LFInst_11_LFInst_2_n19 ,
         \SubCellInst_LFInst_11_LFInst_2_n18 ,
         \SubCellInst_LFInst_11_LFInst_2_n17 ,
         \SubCellInst_LFInst_11_LFInst_2_n16 ,
         \SubCellInst_LFInst_11_LFInst_2_n15 ,
         \SubCellInst_LFInst_11_LFInst_3_n16 ,
         \SubCellInst_LFInst_11_LFInst_3_n15 ,
         \SubCellInst_LFInst_11_LFInst_3_n14 ,
         \SubCellInst_LFInst_11_LFInst_3_n13 ,
         \SubCellInst_LFInst_11_LFInst_3_n12 ,
         \SubCellInst_LFInst_11_LFInst_3_n11 ,
         \SubCellInst_LFInst_12_LFInst_0_n10 ,
         \SubCellInst_LFInst_12_LFInst_0_n9 ,
         \SubCellInst_LFInst_12_LFInst_0_n8 ,
         \SubCellInst_LFInst_12_LFInst_0_n7 ,
         \SubCellInst_LFInst_12_LFInst_1_n18 ,
         \SubCellInst_LFInst_12_LFInst_1_n17 ,
         \SubCellInst_LFInst_12_LFInst_1_n16 ,
         \SubCellInst_LFInst_12_LFInst_1_n15 ,
         \SubCellInst_LFInst_12_LFInst_1_n14 ,
         \SubCellInst_LFInst_12_LFInst_1_n13 ,
         \SubCellInst_LFInst_12_LFInst_1_n12 ,
         \SubCellInst_LFInst_12_LFInst_1_n11 ,
         \SubCellInst_LFInst_12_LFInst_1_n10 ,
         \SubCellInst_LFInst_12_LFInst_2_n22 ,
         \SubCellInst_LFInst_12_LFInst_2_n21 ,
         \SubCellInst_LFInst_12_LFInst_2_n20 ,
         \SubCellInst_LFInst_12_LFInst_2_n19 ,
         \SubCellInst_LFInst_12_LFInst_2_n18 ,
         \SubCellInst_LFInst_12_LFInst_2_n17 ,
         \SubCellInst_LFInst_12_LFInst_2_n16 ,
         \SubCellInst_LFInst_12_LFInst_2_n15 ,
         \SubCellInst_LFInst_12_LFInst_3_n16 ,
         \SubCellInst_LFInst_12_LFInst_3_n15 ,
         \SubCellInst_LFInst_12_LFInst_3_n14 ,
         \SubCellInst_LFInst_12_LFInst_3_n13 ,
         \SubCellInst_LFInst_12_LFInst_3_n12 ,
         \SubCellInst_LFInst_12_LFInst_3_n11 ,
         \SubCellInst_LFInst_13_LFInst_0_n10 ,
         \SubCellInst_LFInst_13_LFInst_0_n9 ,
         \SubCellInst_LFInst_13_LFInst_0_n8 ,
         \SubCellInst_LFInst_13_LFInst_0_n7 ,
         \SubCellInst_LFInst_13_LFInst_1_n18 ,
         \SubCellInst_LFInst_13_LFInst_1_n17 ,
         \SubCellInst_LFInst_13_LFInst_1_n16 ,
         \SubCellInst_LFInst_13_LFInst_1_n15 ,
         \SubCellInst_LFInst_13_LFInst_1_n14 ,
         \SubCellInst_LFInst_13_LFInst_1_n13 ,
         \SubCellInst_LFInst_13_LFInst_1_n12 ,
         \SubCellInst_LFInst_13_LFInst_1_n11 ,
         \SubCellInst_LFInst_13_LFInst_1_n10 ,
         \SubCellInst_LFInst_13_LFInst_2_n22 ,
         \SubCellInst_LFInst_13_LFInst_2_n21 ,
         \SubCellInst_LFInst_13_LFInst_2_n20 ,
         \SubCellInst_LFInst_13_LFInst_2_n19 ,
         \SubCellInst_LFInst_13_LFInst_2_n18 ,
         \SubCellInst_LFInst_13_LFInst_2_n17 ,
         \SubCellInst_LFInst_13_LFInst_2_n16 ,
         \SubCellInst_LFInst_13_LFInst_2_n15 ,
         \SubCellInst_LFInst_13_LFInst_3_n16 ,
         \SubCellInst_LFInst_13_LFInst_3_n15 ,
         \SubCellInst_LFInst_13_LFInst_3_n14 ,
         \SubCellInst_LFInst_13_LFInst_3_n13 ,
         \SubCellInst_LFInst_13_LFInst_3_n12 ,
         \SubCellInst_LFInst_13_LFInst_3_n11 ,
         \SubCellInst_LFInst_14_LFInst_0_n10 ,
         \SubCellInst_LFInst_14_LFInst_0_n9 ,
         \SubCellInst_LFInst_14_LFInst_0_n8 ,
         \SubCellInst_LFInst_14_LFInst_0_n7 ,
         \SubCellInst_LFInst_14_LFInst_1_n18 ,
         \SubCellInst_LFInst_14_LFInst_1_n17 ,
         \SubCellInst_LFInst_14_LFInst_1_n16 ,
         \SubCellInst_LFInst_14_LFInst_1_n15 ,
         \SubCellInst_LFInst_14_LFInst_1_n14 ,
         \SubCellInst_LFInst_14_LFInst_1_n13 ,
         \SubCellInst_LFInst_14_LFInst_1_n12 ,
         \SubCellInst_LFInst_14_LFInst_1_n11 ,
         \SubCellInst_LFInst_14_LFInst_1_n10 ,
         \SubCellInst_LFInst_14_LFInst_2_n22 ,
         \SubCellInst_LFInst_14_LFInst_2_n21 ,
         \SubCellInst_LFInst_14_LFInst_2_n20 ,
         \SubCellInst_LFInst_14_LFInst_2_n19 ,
         \SubCellInst_LFInst_14_LFInst_2_n18 ,
         \SubCellInst_LFInst_14_LFInst_2_n17 ,
         \SubCellInst_LFInst_14_LFInst_2_n16 ,
         \SubCellInst_LFInst_14_LFInst_2_n15 ,
         \SubCellInst_LFInst_14_LFInst_3_n16 ,
         \SubCellInst_LFInst_14_LFInst_3_n15 ,
         \SubCellInst_LFInst_14_LFInst_3_n14 ,
         \SubCellInst_LFInst_14_LFInst_3_n13 ,
         \SubCellInst_LFInst_14_LFInst_3_n12 ,
         \SubCellInst_LFInst_14_LFInst_3_n11 ,
         \SubCellInst_LFInst_15_LFInst_0_n10 ,
         \SubCellInst_LFInst_15_LFInst_0_n9 ,
         \SubCellInst_LFInst_15_LFInst_0_n8 ,
         \SubCellInst_LFInst_15_LFInst_0_n7 ,
         \SubCellInst_LFInst_15_LFInst_1_n18 ,
         \SubCellInst_LFInst_15_LFInst_1_n17 ,
         \SubCellInst_LFInst_15_LFInst_1_n16 ,
         \SubCellInst_LFInst_15_LFInst_1_n15 ,
         \SubCellInst_LFInst_15_LFInst_1_n14 ,
         \SubCellInst_LFInst_15_LFInst_1_n13 ,
         \SubCellInst_LFInst_15_LFInst_1_n12 ,
         \SubCellInst_LFInst_15_LFInst_1_n11 ,
         \SubCellInst_LFInst_15_LFInst_1_n10 ,
         \SubCellInst_LFInst_15_LFInst_2_n22 ,
         \SubCellInst_LFInst_15_LFInst_2_n21 ,
         \SubCellInst_LFInst_15_LFInst_2_n20 ,
         \SubCellInst_LFInst_15_LFInst_2_n19 ,
         \SubCellInst_LFInst_15_LFInst_2_n18 ,
         \SubCellInst_LFInst_15_LFInst_2_n17 ,
         \SubCellInst_LFInst_15_LFInst_2_n16 ,
         \SubCellInst_LFInst_15_LFInst_2_n15 ,
         \SubCellInst_LFInst_15_LFInst_3_n16 ,
         \SubCellInst_LFInst_15_LFInst_3_n15 ,
         \SubCellInst_LFInst_15_LFInst_3_n14 ,
         \SubCellInst_LFInst_15_LFInst_3_n13 ,
         \SubCellInst_LFInst_15_LFInst_3_n12 ,
         \SubCellInst_LFInst_15_LFInst_3_n11 , \MCInst_MC0_v0_2Inst_0_n2 ,
         \MCInst_MC0_v1_2Inst_0_n2 , \MCInst_MC0_v2_3Inst_0_n4 ,
         \MCInst_MC0_v2_3Inst_0_n3 , \MCInst_MC0_v3_3Inst_0_n2 ,
         \MCInst_MC0_v0_2Inst_1_n2 , \MCInst_MC0_v2_1Inst_1_n2 ,
         \MCInst_MC0_v2_2Inst_1_n4 , \MCInst_MC0_v2_2Inst_1_n3 ,
         \MCInst_MC0_v3_3Inst_1_n2 , \MCInst_MC0_v1_1Inst_2_n2 ,
         \MCInst_MC0_v1_2Inst_2_n2 , \MCInst_MC0_v2_1Inst_2_n2 ,
         \MCInst_MC0_v2_2Inst_2_n2 , \MCInst_MC0_v3_1Inst_2_n2 ,
         \MCInst_MC0_v1_2Inst_3_n4 , \MCInst_MC0_v1_2Inst_3_n3 ,
         \MCInst_MC0_v2_2Inst_3_n2 , \MCInst_MC0_v2_3Inst_3_n2 ,
         \MCInst_MC0_r0Inst_XORInst_0_0_n5 ,
         \MCInst_MC0_r0Inst_XORInst_0_0_n4 ,
         \MCInst_MC0_r0Inst_XORInst_0_1_n5 ,
         \MCInst_MC0_r0Inst_XORInst_0_1_n4 ,
         \MCInst_MC0_r0Inst_XORInst_0_2_n5 ,
         \MCInst_MC0_r0Inst_XORInst_0_2_n4 ,
         \MCInst_MC0_r0Inst_XORInst_0_3_n5 ,
         \MCInst_MC0_r0Inst_XORInst_0_3_n4 ,
         \MCInst_MC0_r1Inst_XORInst_0_0_n5 ,
         \MCInst_MC0_r1Inst_XORInst_0_0_n4 ,
         \MCInst_MC0_r1Inst_XORInst_0_1_n5 ,
         \MCInst_MC0_r1Inst_XORInst_0_1_n4 ,
         \MCInst_MC0_r1Inst_XORInst_0_2_n5 ,
         \MCInst_MC0_r1Inst_XORInst_0_2_n4 ,
         \MCInst_MC0_r1Inst_XORInst_0_3_n5 ,
         \MCInst_MC0_r1Inst_XORInst_0_3_n4 ,
         \MCInst_MC0_r2Inst_XORInst_0_0_n5 ,
         \MCInst_MC0_r2Inst_XORInst_0_0_n4 ,
         \MCInst_MC0_r2Inst_XORInst_0_1_n5 ,
         \MCInst_MC0_r2Inst_XORInst_0_1_n4 ,
         \MCInst_MC0_r2Inst_XORInst_0_2_n5 ,
         \MCInst_MC0_r2Inst_XORInst_0_2_n4 ,
         \MCInst_MC0_r2Inst_XORInst_0_3_n5 ,
         \MCInst_MC0_r2Inst_XORInst_0_3_n4 ,
         \MCInst_MC0_r3Inst_XORInst_0_0_n5 ,
         \MCInst_MC0_r3Inst_XORInst_0_0_n4 ,
         \MCInst_MC0_r3Inst_XORInst_0_1_n5 ,
         \MCInst_MC0_r3Inst_XORInst_0_1_n4 ,
         \MCInst_MC0_r3Inst_XORInst_0_2_n5 ,
         \MCInst_MC0_r3Inst_XORInst_0_2_n4 ,
         \MCInst_MC0_r3Inst_XORInst_0_3_n5 ,
         \MCInst_MC0_r3Inst_XORInst_0_3_n4 , \MCInst_MC1_v0_2Inst_0_n2 ,
         \MCInst_MC1_v1_2Inst_0_n2 , \MCInst_MC1_v2_3Inst_0_n4 ,
         \MCInst_MC1_v2_3Inst_0_n3 , \MCInst_MC1_v3_3Inst_0_n2 ,
         \MCInst_MC1_v0_2Inst_1_n2 , \MCInst_MC1_v2_1Inst_1_n2 ,
         \MCInst_MC1_v2_2Inst_1_n4 , \MCInst_MC1_v2_2Inst_1_n3 ,
         \MCInst_MC1_v3_3Inst_1_n2 , \MCInst_MC1_v1_1Inst_2_n2 ,
         \MCInst_MC1_v1_2Inst_2_n2 , \MCInst_MC1_v2_1Inst_2_n2 ,
         \MCInst_MC1_v2_2Inst_2_n2 , \MCInst_MC1_v3_1Inst_2_n2 ,
         \MCInst_MC1_v1_2Inst_3_n4 , \MCInst_MC1_v1_2Inst_3_n3 ,
         \MCInst_MC1_v2_2Inst_3_n2 , \MCInst_MC1_v2_3Inst_3_n2 ,
         \MCInst_MC1_r0Inst_XORInst_0_0_n5 ,
         \MCInst_MC1_r0Inst_XORInst_0_0_n4 ,
         \MCInst_MC1_r0Inst_XORInst_0_1_n5 ,
         \MCInst_MC1_r0Inst_XORInst_0_1_n4 ,
         \MCInst_MC1_r0Inst_XORInst_0_2_n5 ,
         \MCInst_MC1_r0Inst_XORInst_0_2_n4 ,
         \MCInst_MC1_r0Inst_XORInst_0_3_n5 ,
         \MCInst_MC1_r0Inst_XORInst_0_3_n4 ,
         \MCInst_MC1_r1Inst_XORInst_0_0_n5 ,
         \MCInst_MC1_r1Inst_XORInst_0_0_n4 ,
         \MCInst_MC1_r1Inst_XORInst_0_1_n5 ,
         \MCInst_MC1_r1Inst_XORInst_0_1_n4 ,
         \MCInst_MC1_r1Inst_XORInst_0_2_n5 ,
         \MCInst_MC1_r1Inst_XORInst_0_2_n4 ,
         \MCInst_MC1_r1Inst_XORInst_0_3_n5 ,
         \MCInst_MC1_r1Inst_XORInst_0_3_n4 ,
         \MCInst_MC1_r2Inst_XORInst_0_0_n5 ,
         \MCInst_MC1_r2Inst_XORInst_0_0_n4 ,
         \MCInst_MC1_r2Inst_XORInst_0_1_n5 ,
         \MCInst_MC1_r2Inst_XORInst_0_1_n4 ,
         \MCInst_MC1_r2Inst_XORInst_0_2_n5 ,
         \MCInst_MC1_r2Inst_XORInst_0_2_n4 ,
         \MCInst_MC1_r2Inst_XORInst_0_3_n5 ,
         \MCInst_MC1_r2Inst_XORInst_0_3_n4 ,
         \MCInst_MC1_r3Inst_XORInst_0_0_n5 ,
         \MCInst_MC1_r3Inst_XORInst_0_0_n4 ,
         \MCInst_MC1_r3Inst_XORInst_0_1_n5 ,
         \MCInst_MC1_r3Inst_XORInst_0_1_n4 ,
         \MCInst_MC1_r3Inst_XORInst_0_2_n5 ,
         \MCInst_MC1_r3Inst_XORInst_0_2_n4 ,
         \MCInst_MC1_r3Inst_XORInst_0_3_n5 ,
         \MCInst_MC1_r3Inst_XORInst_0_3_n4 , \MCInst_MC2_v0_2Inst_0_n2 ,
         \MCInst_MC2_v1_2Inst_0_n2 , \MCInst_MC2_v2_3Inst_0_n4 ,
         \MCInst_MC2_v2_3Inst_0_n3 , \MCInst_MC2_v3_3Inst_0_n2 ,
         \MCInst_MC2_v0_2Inst_1_n2 , \MCInst_MC2_v2_1Inst_1_n2 ,
         \MCInst_MC2_v2_2Inst_1_n4 , \MCInst_MC2_v2_2Inst_1_n3 ,
         \MCInst_MC2_v3_3Inst_1_n2 , \MCInst_MC2_v1_1Inst_2_n2 ,
         \MCInst_MC2_v1_2Inst_2_n2 , \MCInst_MC2_v2_1Inst_2_n2 ,
         \MCInst_MC2_v2_2Inst_2_n2 , \MCInst_MC2_v3_1Inst_2_n2 ,
         \MCInst_MC2_v1_2Inst_3_n4 , \MCInst_MC2_v1_2Inst_3_n3 ,
         \MCInst_MC2_v2_2Inst_3_n2 , \MCInst_MC2_v2_3Inst_3_n2 ,
         \MCInst_MC2_r0Inst_XORInst_0_0_n5 ,
         \MCInst_MC2_r0Inst_XORInst_0_0_n4 ,
         \MCInst_MC2_r0Inst_XORInst_0_1_n5 ,
         \MCInst_MC2_r0Inst_XORInst_0_1_n4 ,
         \MCInst_MC2_r0Inst_XORInst_0_2_n5 ,
         \MCInst_MC2_r0Inst_XORInst_0_2_n4 ,
         \MCInst_MC2_r0Inst_XORInst_0_3_n5 ,
         \MCInst_MC2_r0Inst_XORInst_0_3_n4 ,
         \MCInst_MC2_r1Inst_XORInst_0_0_n5 ,
         \MCInst_MC2_r1Inst_XORInst_0_0_n4 ,
         \MCInst_MC2_r1Inst_XORInst_0_1_n5 ,
         \MCInst_MC2_r1Inst_XORInst_0_1_n4 ,
         \MCInst_MC2_r1Inst_XORInst_0_2_n5 ,
         \MCInst_MC2_r1Inst_XORInst_0_2_n4 ,
         \MCInst_MC2_r1Inst_XORInst_0_3_n5 ,
         \MCInst_MC2_r1Inst_XORInst_0_3_n4 ,
         \MCInst_MC2_r2Inst_XORInst_0_0_n5 ,
         \MCInst_MC2_r2Inst_XORInst_0_0_n4 ,
         \MCInst_MC2_r2Inst_XORInst_0_1_n5 ,
         \MCInst_MC2_r2Inst_XORInst_0_1_n4 ,
         \MCInst_MC2_r2Inst_XORInst_0_2_n5 ,
         \MCInst_MC2_r2Inst_XORInst_0_2_n4 ,
         \MCInst_MC2_r2Inst_XORInst_0_3_n5 ,
         \MCInst_MC2_r2Inst_XORInst_0_3_n4 ,
         \MCInst_MC2_r3Inst_XORInst_0_0_n5 ,
         \MCInst_MC2_r3Inst_XORInst_0_0_n4 ,
         \MCInst_MC2_r3Inst_XORInst_0_1_n5 ,
         \MCInst_MC2_r3Inst_XORInst_0_1_n4 ,
         \MCInst_MC2_r3Inst_XORInst_0_2_n5 ,
         \MCInst_MC2_r3Inst_XORInst_0_2_n4 ,
         \MCInst_MC2_r3Inst_XORInst_0_3_n5 ,
         \MCInst_MC2_r3Inst_XORInst_0_3_n4 , \MCInst_MC3_v0_2Inst_0_n2 ,
         \MCInst_MC3_v1_2Inst_0_n2 , \MCInst_MC3_v2_3Inst_0_n4 ,
         \MCInst_MC3_v2_3Inst_0_n3 , \MCInst_MC3_v3_3Inst_0_n2 ,
         \MCInst_MC3_v0_2Inst_1_n2 , \MCInst_MC3_v2_1Inst_1_n2 ,
         \MCInst_MC3_v2_2Inst_1_n4 , \MCInst_MC3_v2_2Inst_1_n3 ,
         \MCInst_MC3_v3_3Inst_1_n2 , \MCInst_MC3_v1_1Inst_2_n2 ,
         \MCInst_MC3_v1_2Inst_2_n2 , \MCInst_MC3_v2_1Inst_2_n2 ,
         \MCInst_MC3_v2_2Inst_2_n2 , \MCInst_MC3_v3_1Inst_2_n2 ,
         \MCInst_MC3_v1_2Inst_3_n4 , \MCInst_MC3_v1_2Inst_3_n3 ,
         \MCInst_MC3_v2_2Inst_3_n2 , \MCInst_MC3_v2_3Inst_3_n2 ,
         \MCInst_MC3_r0Inst_XORInst_0_0_n5 ,
         \MCInst_MC3_r0Inst_XORInst_0_0_n4 ,
         \MCInst_MC3_r0Inst_XORInst_0_1_n5 ,
         \MCInst_MC3_r0Inst_XORInst_0_1_n4 ,
         \MCInst_MC3_r0Inst_XORInst_0_2_n5 ,
         \MCInst_MC3_r0Inst_XORInst_0_2_n4 ,
         \MCInst_MC3_r0Inst_XORInst_0_3_n5 ,
         \MCInst_MC3_r0Inst_XORInst_0_3_n4 ,
         \MCInst_MC3_r1Inst_XORInst_0_0_n5 ,
         \MCInst_MC3_r1Inst_XORInst_0_0_n4 ,
         \MCInst_MC3_r1Inst_XORInst_0_1_n5 ,
         \MCInst_MC3_r1Inst_XORInst_0_1_n4 ,
         \MCInst_MC3_r1Inst_XORInst_0_2_n5 ,
         \MCInst_MC3_r1Inst_XORInst_0_2_n4 ,
         \MCInst_MC3_r1Inst_XORInst_0_3_n5 ,
         \MCInst_MC3_r1Inst_XORInst_0_3_n4 ,
         \MCInst_MC3_r2Inst_XORInst_0_0_n5 ,
         \MCInst_MC3_r2Inst_XORInst_0_0_n4 ,
         \MCInst_MC3_r2Inst_XORInst_0_1_n5 ,
         \MCInst_MC3_r2Inst_XORInst_0_1_n4 ,
         \MCInst_MC3_r2Inst_XORInst_0_2_n5 ,
         \MCInst_MC3_r2Inst_XORInst_0_2_n4 ,
         \MCInst_MC3_r2Inst_XORInst_0_3_n5 ,
         \MCInst_MC3_r2Inst_XORInst_0_3_n4 ,
         \MCInst_MC3_r3Inst_XORInst_0_0_n5 ,
         \MCInst_MC3_r3Inst_XORInst_0_0_n4 ,
         \MCInst_MC3_r3Inst_XORInst_0_1_n5 ,
         \MCInst_MC3_r3Inst_XORInst_0_1_n4 ,
         \MCInst_MC3_r3Inst_XORInst_0_2_n5 ,
         \MCInst_MC3_r3Inst_XORInst_0_2_n4 ,
         \MCInst_MC3_r3Inst_XORInst_0_3_n5 ,
         \MCInst_MC3_r3Inst_XORInst_0_3_n4 ,
         \Red_PlaintextInst_LFInst_0_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_0_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_0_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_1_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_1_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_1_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_2_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_2_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_2_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_3_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_3_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_3_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_4_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_4_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_4_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_5_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_5_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_5_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_6_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_6_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_6_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_7_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_7_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_7_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_8_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_8_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_8_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_9_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_9_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_9_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_10_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_10_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_10_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_11_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_11_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_11_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_12_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_12_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_12_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_13_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_13_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_13_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_14_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_14_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_14_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_15_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_15_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_15_LFInst_2_n2 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n7 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n6 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n5 ,
         \Red_SubCellInst_LFInst_0_LFInst_1_n4 ,
         \Red_SubCellInst_LFInst_0_LFInst_1_n3 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n11 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n10 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n9 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n8 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n7 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n7 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n6 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n5 ,
         \Red_SubCellInst_LFInst_1_LFInst_1_n4 ,
         \Red_SubCellInst_LFInst_1_LFInst_1_n3 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n11 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n10 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n9 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n8 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n7 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n7 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n6 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n5 ,
         \Red_SubCellInst_LFInst_2_LFInst_1_n4 ,
         \Red_SubCellInst_LFInst_2_LFInst_1_n3 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n11 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n10 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n9 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n8 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n7 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n7 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n6 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n5 ,
         \Red_SubCellInst_LFInst_3_LFInst_1_n4 ,
         \Red_SubCellInst_LFInst_3_LFInst_1_n3 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n11 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n10 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n9 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n8 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n7 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n7 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n6 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n5 ,
         \Red_SubCellInst_LFInst_4_LFInst_1_n4 ,
         \Red_SubCellInst_LFInst_4_LFInst_1_n3 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n11 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n10 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n9 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n8 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n7 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n7 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n6 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n5 ,
         \Red_SubCellInst_LFInst_5_LFInst_1_n4 ,
         \Red_SubCellInst_LFInst_5_LFInst_1_n3 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n11 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n10 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n9 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n8 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n7 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n7 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n6 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n5 ,
         \Red_SubCellInst_LFInst_6_LFInst_1_n4 ,
         \Red_SubCellInst_LFInst_6_LFInst_1_n3 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n11 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n10 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n9 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n8 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n7 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n7 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n6 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n5 ,
         \Red_SubCellInst_LFInst_7_LFInst_1_n4 ,
         \Red_SubCellInst_LFInst_7_LFInst_1_n3 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n11 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n10 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n9 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n8 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n7 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n7 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n6 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n5 ,
         \Red_SubCellInst_LFInst_8_LFInst_1_n4 ,
         \Red_SubCellInst_LFInst_8_LFInst_1_n3 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n11 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n10 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n9 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n8 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n7 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n7 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n6 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n5 ,
         \Red_SubCellInst_LFInst_9_LFInst_1_n4 ,
         \Red_SubCellInst_LFInst_9_LFInst_1_n3 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n11 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n10 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n9 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n8 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n7 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n7 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n6 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n5 ,
         \Red_SubCellInst_LFInst_10_LFInst_1_n4 ,
         \Red_SubCellInst_LFInst_10_LFInst_1_n3 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n11 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n10 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n9 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n8 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n7 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n7 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n6 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n5 ,
         \Red_SubCellInst_LFInst_11_LFInst_1_n4 ,
         \Red_SubCellInst_LFInst_11_LFInst_1_n3 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n11 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n10 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n9 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n8 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n7 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n7 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n6 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n5 ,
         \Red_SubCellInst_LFInst_12_LFInst_1_n4 ,
         \Red_SubCellInst_LFInst_12_LFInst_1_n3 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n11 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n10 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n9 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n8 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n7 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n7 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n6 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n5 ,
         \Red_SubCellInst_LFInst_13_LFInst_1_n4 ,
         \Red_SubCellInst_LFInst_13_LFInst_1_n3 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n11 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n10 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n9 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n8 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n7 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n7 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n6 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n5 ,
         \Red_SubCellInst_LFInst_14_LFInst_1_n4 ,
         \Red_SubCellInst_LFInst_14_LFInst_1_n3 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n11 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n10 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n9 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n8 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n7 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n7 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n6 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n5 ,
         \Red_SubCellInst_LFInst_15_LFInst_1_n4 ,
         \Red_SubCellInst_LFInst_15_LFInst_1_n3 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n11 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n10 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n9 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n8 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n7 ,
         \Red_MCInst_MC0_v1_0Inst_0_n2 , \Red_MCInst_MC0_v2_2Inst_0_n2 ,
         \Red_MCInst_MC0_v2_3Inst_0_n2 , \Red_MCInst_MC0_v3_2Inst_0_n4 ,
         \Red_MCInst_MC0_v3_2Inst_0_n3 , \Red_MCInst_MC0_v0_1Inst_1_n2 ,
         \Red_MCInst_MC0_v1_0Inst_1_n2 , \Red_MCInst_MC0_v1_1Inst_1_n4 ,
         \Red_MCInst_MC0_v1_1Inst_1_n3 , \Red_MCInst_MC0_v3_1Inst_1_n4 ,
         \Red_MCInst_MC0_v3_1Inst_1_n3 , \Red_MCInst_MC0_v0_0Inst_2_n2 ,
         \Red_MCInst_MC0_v0_3Inst_2_n4 , \Red_MCInst_MC0_v0_3Inst_2_n3 ,
         \Red_MCInst_MC0_v1_0Inst_2_n2 , \Red_MCInst_MC0_v1_2Inst_2_n2 ,
         \Red_MCInst_MC0_v1_3Inst_2_n4 , \Red_MCInst_MC0_v1_3Inst_2_n3 ,
         \Red_MCInst_MC0_v2_0Inst_2_n4 , \Red_MCInst_MC0_v2_0Inst_2_n3 ,
         \Red_MCInst_MC0_v3_0Inst_2_n4 , \Red_MCInst_MC0_v3_0Inst_2_n3 ,
         \Red_MCInst_MC0_v3_2Inst_2_n2 ,
         \Red_MCInst_MC0_r0Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC0_r0Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC0_r0Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC0_r0Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC0_r0Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC0_r0Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC0_r1Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC0_r1Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC0_r1Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC0_r1Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC0_r1Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC0_r1Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC0_r2Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC0_r2Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC0_r2Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC0_r2Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC0_r2Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC0_r2Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC0_r3Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC0_r3Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC0_r3Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC0_r3Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC0_r3Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC0_r3Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC1_v1_0Inst_0_n2 , \Red_MCInst_MC1_v2_2Inst_0_n2 ,
         \Red_MCInst_MC1_v2_3Inst_0_n2 , \Red_MCInst_MC1_v3_2Inst_0_n4 ,
         \Red_MCInst_MC1_v3_2Inst_0_n3 , \Red_MCInst_MC1_v0_1Inst_1_n2 ,
         \Red_MCInst_MC1_v1_0Inst_1_n2 , \Red_MCInst_MC1_v1_1Inst_1_n4 ,
         \Red_MCInst_MC1_v1_1Inst_1_n3 , \Red_MCInst_MC1_v3_1Inst_1_n4 ,
         \Red_MCInst_MC1_v3_1Inst_1_n3 , \Red_MCInst_MC1_v0_0Inst_2_n2 ,
         \Red_MCInst_MC1_v0_3Inst_2_n4 , \Red_MCInst_MC1_v0_3Inst_2_n3 ,
         \Red_MCInst_MC1_v1_0Inst_2_n2 , \Red_MCInst_MC1_v1_2Inst_2_n2 ,
         \Red_MCInst_MC1_v1_3Inst_2_n4 , \Red_MCInst_MC1_v1_3Inst_2_n3 ,
         \Red_MCInst_MC1_v2_0Inst_2_n4 , \Red_MCInst_MC1_v2_0Inst_2_n3 ,
         \Red_MCInst_MC1_v3_0Inst_2_n4 , \Red_MCInst_MC1_v3_0Inst_2_n3 ,
         \Red_MCInst_MC1_v3_2Inst_2_n2 ,
         \Red_MCInst_MC1_r0Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC1_r0Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC1_r0Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC1_r0Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC1_r0Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC1_r0Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC1_r1Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC1_r1Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC1_r1Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC1_r1Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC1_r1Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC1_r1Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC1_r2Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC1_r2Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC1_r2Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC1_r2Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC1_r2Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC1_r2Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC1_r3Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC1_r3Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC1_r3Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC1_r3Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC1_r3Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC1_r3Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC2_v1_0Inst_0_n2 , \Red_MCInst_MC2_v2_2Inst_0_n2 ,
         \Red_MCInst_MC2_v2_3Inst_0_n2 , \Red_MCInst_MC2_v3_2Inst_0_n4 ,
         \Red_MCInst_MC2_v3_2Inst_0_n3 , \Red_MCInst_MC2_v0_1Inst_1_n2 ,
         \Red_MCInst_MC2_v1_0Inst_1_n2 , \Red_MCInst_MC2_v1_1Inst_1_n4 ,
         \Red_MCInst_MC2_v1_1Inst_1_n3 , \Red_MCInst_MC2_v3_1Inst_1_n4 ,
         \Red_MCInst_MC2_v3_1Inst_1_n3 , \Red_MCInst_MC2_v0_0Inst_2_n2 ,
         \Red_MCInst_MC2_v0_3Inst_2_n4 , \Red_MCInst_MC2_v0_3Inst_2_n3 ,
         \Red_MCInst_MC2_v1_0Inst_2_n2 , \Red_MCInst_MC2_v1_2Inst_2_n2 ,
         \Red_MCInst_MC2_v1_3Inst_2_n4 , \Red_MCInst_MC2_v1_3Inst_2_n3 ,
         \Red_MCInst_MC2_v2_0Inst_2_n4 , \Red_MCInst_MC2_v2_0Inst_2_n3 ,
         \Red_MCInst_MC2_v3_0Inst_2_n4 , \Red_MCInst_MC2_v3_0Inst_2_n3 ,
         \Red_MCInst_MC2_v3_2Inst_2_n2 ,
         \Red_MCInst_MC2_r0Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC2_r0Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC2_r0Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC2_r0Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC2_r0Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC2_r0Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC2_r1Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC2_r1Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC2_r1Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC2_r1Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC2_r1Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC2_r1Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC2_r2Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC2_r2Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC2_r2Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC2_r2Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC2_r2Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC2_r2Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC2_r3Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC2_r3Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC2_r3Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC2_r3Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC2_r3Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC2_r3Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC3_v1_0Inst_0_n2 , \Red_MCInst_MC3_v2_2Inst_0_n2 ,
         \Red_MCInst_MC3_v2_3Inst_0_n2 , \Red_MCInst_MC3_v3_2Inst_0_n4 ,
         \Red_MCInst_MC3_v3_2Inst_0_n3 , \Red_MCInst_MC3_v0_1Inst_1_n2 ,
         \Red_MCInst_MC3_v1_0Inst_1_n2 , \Red_MCInst_MC3_v1_1Inst_1_n4 ,
         \Red_MCInst_MC3_v1_1Inst_1_n3 , \Red_MCInst_MC3_v3_1Inst_1_n4 ,
         \Red_MCInst_MC3_v3_1Inst_1_n3 , \Red_MCInst_MC3_v0_0Inst_2_n2 ,
         \Red_MCInst_MC3_v0_3Inst_2_n4 , \Red_MCInst_MC3_v0_3Inst_2_n3 ,
         \Red_MCInst_MC3_v1_0Inst_2_n2 , \Red_MCInst_MC3_v1_2Inst_2_n2 ,
         \Red_MCInst_MC3_v1_3Inst_2_n4 , \Red_MCInst_MC3_v1_3Inst_2_n3 ,
         \Red_MCInst_MC3_v2_0Inst_2_n4 , \Red_MCInst_MC3_v2_0Inst_2_n3 ,
         \Red_MCInst_MC3_v3_0Inst_2_n4 , \Red_MCInst_MC3_v3_0Inst_2_n3 ,
         \Red_MCInst_MC3_v3_2Inst_2_n2 ,
         \Red_MCInst_MC3_r0Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC3_r0Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC3_r0Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC3_r0Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC3_r0Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC3_r0Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC3_r1Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC3_r1Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC3_r1Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC3_r1Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC3_r1Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC3_r1Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC3_r2Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC3_r2Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC3_r2Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC3_r2Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC3_r2Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC3_r2Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC3_r3Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC3_r3Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC3_r3Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC3_r3Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC3_r3Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC3_r3Inst_XORInst_0_2_n4 ,
         \Red_ToCheckInst_LFInst_0_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_0_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_0_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_1_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_1_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_1_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_2_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_2_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_2_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_3_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_3_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_3_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_4_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_4_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_4_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_5_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_5_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_5_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_6_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_6_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_6_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_7_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_7_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_7_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_8_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_8_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_8_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_9_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_9_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_9_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_10_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_10_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_10_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_11_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_11_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_11_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_12_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_12_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_12_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_13_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_13_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_13_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_14_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_14_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_14_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_15_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_15_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_15_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_16_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_16_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_16_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_17_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_17_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_17_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_18_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_18_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_18_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_19_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_19_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_19_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_20_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_20_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_20_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_21_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_21_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_21_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_22_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_22_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_22_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_23_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_23_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_23_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_24_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_24_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_24_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_25_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_25_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_25_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_26_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_26_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_26_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_27_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_27_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_27_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_28_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_28_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_28_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_29_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_29_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_29_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_30_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_30_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_30_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_31_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_31_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_31_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_32_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_32_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_32_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_33_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_33_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_33_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_34_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_34_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_34_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_35_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_35_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_35_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_36_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_36_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_36_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_37_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_37_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_37_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_38_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_38_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_38_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_39_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_39_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_39_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_40_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_40_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_40_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_41_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_41_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_41_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_42_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_42_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_42_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_43_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_43_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_43_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_44_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_44_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_44_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_45_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_45_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_45_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_46_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_46_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_46_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_47_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_47_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_47_LFInst_2_n2 , \Check1_CheckInst_0_n94 ,
         \Check1_CheckInst_0_n93 , \Check1_CheckInst_0_n92 ,
         \Check1_CheckInst_0_n91 , \Check1_CheckInst_0_n90 ,
         \Check1_CheckInst_0_n89 , \Check1_CheckInst_0_n88 ,
         \Check1_CheckInst_0_n87 , \Check1_CheckInst_0_n86 ,
         \Check1_CheckInst_0_n85 , \Check1_CheckInst_0_n84 ,
         \Check1_CheckInst_0_n83 , \Check1_CheckInst_0_n82 ,
         \Check1_CheckInst_0_n81 , \Check1_CheckInst_0_n80 ,
         \Check1_CheckInst_0_n79 , \Check1_CheckInst_0_n78 ,
         \Check1_CheckInst_0_n77 , \Check1_CheckInst_0_n76 ,
         \Check1_CheckInst_0_n75 , \Check1_CheckInst_0_n74 ,
         \Check1_CheckInst_0_n73 , \Check1_CheckInst_0_n72 ,
         \Check1_CheckInst_0_n71 , \Check1_CheckInst_0_n70 ,
         \Check1_CheckInst_0_n69 , \Check1_CheckInst_0_n68 ,
         \Check1_CheckInst_0_n67 , \Check1_CheckInst_0_n66 ,
         \Check1_CheckInst_0_n65 , \Check1_CheckInst_0_n64 ,
         \Check1_CheckInst_0_n63 , \Check1_CheckInst_0_n62 ,
         \Check1_CheckInst_0_n61 , \Check1_CheckInst_0_n60 ,
         \Check1_CheckInst_0_n59 , \Check1_CheckInst_0_n58 ,
         \Check1_CheckInst_0_n57 , \Check1_CheckInst_0_n56 ,
         \Check1_CheckInst_0_n55 , \Check1_CheckInst_0_n54 ,
         \Check1_CheckInst_0_n53 , \Check1_CheckInst_0_n52 ,
         \Check1_CheckInst_0_n51 , \Check1_CheckInst_0_n50 ,
         \Check1_CheckInst_0_n49 , \Check1_CheckInst_0_n48 ,
         \Check1_CheckInst_0_n47 , \Check1_CheckInst_0_n46 ,
         \Check1_CheckInst_0_n45 , \Check1_CheckInst_0_n44 ,
         \Check1_CheckInst_0_n43 , \Check1_CheckInst_0_n42 ,
         \Check1_CheckInst_0_n41 , \Check1_CheckInst_0_n40 ,
         \Check1_CheckInst_0_n39 , \Check1_CheckInst_0_n38 ,
         \Check1_CheckInst_0_n37 , \Check1_CheckInst_0_n36 ,
         \Check1_CheckInst_0_n35 , \Check1_CheckInst_0_n34 ,
         \Check1_CheckInst_0_n33 , \Check1_CheckInst_0_n32 ,
         \Check1_CheckInst_0_n31 , \Check1_CheckInst_0_n30 ,
         \Check1_CheckInst_0_n29 , \Check1_CheckInst_0_n28 ,
         \Check1_CheckInst_0_n27 , \Check1_CheckInst_0_n26 ,
         \Check1_CheckInst_0_n25 , \Check1_CheckInst_0_n24 ,
         \Check1_CheckInst_0_n23 , \Check1_CheckInst_0_n22 ,
         \Check1_CheckInst_0_n21 , \Check1_CheckInst_0_n20 ,
         \Check1_CheckInst_0_n19 , \Check1_CheckInst_0_n18 ,
         \Check1_CheckInst_0_n17 , \Check1_CheckInst_0_n16 ,
         \Check1_CheckInst_0_n15 , \Check1_CheckInst_0_n14 ,
         \Check1_CheckInst_0_n13 , \Check1_CheckInst_0_n12 ,
         \Check1_CheckInst_0_n11 , \Check1_CheckInst_0_n10 ,
         \Check1_CheckInst_0_n9 , \Check1_CheckInst_0_n8 ,
         \Check1_CheckInst_0_n7 , \Check1_CheckInst_0_n6 ,
         \Check1_CheckInst_0_n5 , \Check1_CheckInst_0_n4 ,
         \Check1_CheckInst_0_n3 , \Check1_CheckInst_0_n2 ,
         \Check1_CheckInst_0_n1 , \Check1_CheckInst_1_n96 ,
         \Check1_CheckInst_1_n95 , \Check1_CheckInst_1_n94 ,
         \Check1_CheckInst_1_n93 , \Check1_CheckInst_1_n92 ,
         \Check1_CheckInst_1_n91 , \Check1_CheckInst_1_n90 ,
         \Check1_CheckInst_1_n89 , \Check1_CheckInst_1_n88 ,
         \Check1_CheckInst_1_n87 , \Check1_CheckInst_1_n86 ,
         \Check1_CheckInst_1_n85 , \Check1_CheckInst_1_n84 ,
         \Check1_CheckInst_1_n83 , \Check1_CheckInst_1_n82 ,
         \Check1_CheckInst_1_n81 , \Check1_CheckInst_1_n80 ,
         \Check1_CheckInst_1_n79 , \Check1_CheckInst_1_n78 ,
         \Check1_CheckInst_1_n77 , \Check1_CheckInst_1_n76 ,
         \Check1_CheckInst_1_n75 , \Check1_CheckInst_1_n74 ,
         \Check1_CheckInst_1_n73 , \Check1_CheckInst_1_n72 ,
         \Check1_CheckInst_1_n71 , \Check1_CheckInst_1_n70 ,
         \Check1_CheckInst_1_n69 , \Check1_CheckInst_1_n68 ,
         \Check1_CheckInst_1_n67 , \Check1_CheckInst_1_n66 ,
         \Check1_CheckInst_1_n65 , \Check1_CheckInst_1_n64 ,
         \Check1_CheckInst_1_n63 , \Check1_CheckInst_1_n62 ,
         \Check1_CheckInst_1_n61 , \Check1_CheckInst_1_n60 ,
         \Check1_CheckInst_1_n59 , \Check1_CheckInst_1_n58 ,
         \Check1_CheckInst_1_n57 , \Check1_CheckInst_1_n56 ,
         \Check1_CheckInst_1_n55 , \Check1_CheckInst_1_n54 ,
         \Check1_CheckInst_1_n53 , \Check1_CheckInst_1_n52 ,
         \Check1_CheckInst_1_n51 , \Check1_CheckInst_1_n50 ,
         \Check1_CheckInst_1_n49 , \Check1_CheckInst_1_n48 ,
         \Check1_CheckInst_1_n47 , \Check1_CheckInst_1_n46 ,
         \Check1_CheckInst_1_n45 , \Check1_CheckInst_1_n44 ,
         \Check1_CheckInst_1_n43 , \Check1_CheckInst_1_n42 ,
         \Check1_CheckInst_1_n41 , \Check1_CheckInst_1_n40 ,
         \Check1_CheckInst_1_n39 , \Check1_CheckInst_1_n38 ,
         \Check1_CheckInst_1_n37 , \Check1_CheckInst_1_n36 ,
         \Check1_CheckInst_1_n35 , \Check1_CheckInst_1_n34 ,
         \Check1_CheckInst_1_n33 , \Check1_CheckInst_1_n32 ,
         \Check1_CheckInst_1_n31 , \Check1_CheckInst_1_n30 ,
         \Check1_CheckInst_1_n29 , \Check1_CheckInst_1_n28 ,
         \Check1_CheckInst_1_n27 , \Check1_CheckInst_1_n26 ,
         \Check1_CheckInst_1_n25 , \Check1_CheckInst_1_n24 ,
         \Check1_CheckInst_1_n23 , \Check1_CheckInst_1_n22 ,
         \Check1_CheckInst_1_n21 , \Check1_CheckInst_1_n20 ,
         \Check1_CheckInst_1_n19 , \Check1_CheckInst_1_n18 ,
         \Check1_CheckInst_1_n17 , \Check1_CheckInst_1_n16 ,
         \Check1_CheckInst_1_n15 , \Check1_CheckInst_1_n14 ,
         \Check1_CheckInst_1_n13 , \Check1_CheckInst_1_n12 ,
         \Check1_CheckInst_1_n11 , \Check1_CheckInst_1_n10 ,
         \Check1_CheckInst_1_n9 , \Check1_CheckInst_1_n8 ,
         \Check1_CheckInst_1_n7 , \Check1_CheckInst_1_n6 ,
         \Check1_CheckInst_1_n5 , \Check1_CheckInst_1_n4 ,
         \Check1_CheckInst_1_n3 , \Check1_CheckInst_2_n96 ,
         \Check1_CheckInst_2_n95 , \Check1_CheckInst_2_n94 ,
         \Check1_CheckInst_2_n93 , \Check1_CheckInst_2_n92 ,
         \Check1_CheckInst_2_n91 , \Check1_CheckInst_2_n90 ,
         \Check1_CheckInst_2_n89 , \Check1_CheckInst_2_n88 ,
         \Check1_CheckInst_2_n87 , \Check1_CheckInst_2_n86 ,
         \Check1_CheckInst_2_n85 , \Check1_CheckInst_2_n84 ,
         \Check1_CheckInst_2_n83 , \Check1_CheckInst_2_n82 ,
         \Check1_CheckInst_2_n81 , \Check1_CheckInst_2_n80 ,
         \Check1_CheckInst_2_n79 , \Check1_CheckInst_2_n78 ,
         \Check1_CheckInst_2_n77 , \Check1_CheckInst_2_n76 ,
         \Check1_CheckInst_2_n75 , \Check1_CheckInst_2_n74 ,
         \Check1_CheckInst_2_n73 , \Check1_CheckInst_2_n72 ,
         \Check1_CheckInst_2_n71 , \Check1_CheckInst_2_n70 ,
         \Check1_CheckInst_2_n69 , \Check1_CheckInst_2_n68 ,
         \Check1_CheckInst_2_n67 , \Check1_CheckInst_2_n66 ,
         \Check1_CheckInst_2_n65 , \Check1_CheckInst_2_n64 ,
         \Check1_CheckInst_2_n63 , \Check1_CheckInst_2_n62 ,
         \Check1_CheckInst_2_n61 , \Check1_CheckInst_2_n60 ,
         \Check1_CheckInst_2_n59 , \Check1_CheckInst_2_n58 ,
         \Check1_CheckInst_2_n57 , \Check1_CheckInst_2_n56 ,
         \Check1_CheckInst_2_n55 , \Check1_CheckInst_2_n54 ,
         \Check1_CheckInst_2_n53 , \Check1_CheckInst_2_n52 ,
         \Check1_CheckInst_2_n51 , \Check1_CheckInst_2_n50 ,
         \Check1_CheckInst_2_n49 , \Check1_CheckInst_2_n48 ,
         \Check1_CheckInst_2_n47 , \Check1_CheckInst_2_n46 ,
         \Check1_CheckInst_2_n45 , \Check1_CheckInst_2_n44 ,
         \Check1_CheckInst_2_n43 , \Check1_CheckInst_2_n42 ,
         \Check1_CheckInst_2_n41 , \Check1_CheckInst_2_n40 ,
         \Check1_CheckInst_2_n39 , \Check1_CheckInst_2_n38 ,
         \Check1_CheckInst_2_n37 , \Check1_CheckInst_2_n36 ,
         \Check1_CheckInst_2_n35 , \Check1_CheckInst_2_n34 ,
         \Check1_CheckInst_2_n33 , \Check1_CheckInst_2_n32 ,
         \Check1_CheckInst_2_n31 , \Check1_CheckInst_2_n30 ,
         \Check1_CheckInst_2_n29 , \Check1_CheckInst_2_n28 ,
         \Check1_CheckInst_2_n27 , \Check1_CheckInst_2_n26 ,
         \Check1_CheckInst_2_n25 , \Check1_CheckInst_2_n24 ,
         \Check1_CheckInst_2_n23 , \Check1_CheckInst_2_n22 ,
         \Check1_CheckInst_2_n21 , \Check1_CheckInst_2_n20 ,
         \Check1_CheckInst_2_n19 , \Check1_CheckInst_2_n18 ,
         \Check1_CheckInst_2_n17 , \Check1_CheckInst_2_n16 ,
         \Check1_CheckInst_2_n15 , \Check1_CheckInst_2_n14 ,
         \Check1_CheckInst_2_n13 , \Check1_CheckInst_2_n12 ,
         \Check1_CheckInst_2_n11 , \Check1_CheckInst_2_n10 ,
         \Check1_CheckInst_2_n9 , \Check1_CheckInst_2_n8 ,
         \Check1_CheckInst_2_n7 , \Check1_CheckInst_2_n6 ,
         \Check1_CheckInst_2_n5 , \Check1_CheckInst_2_n4 ,
         \Check1_CheckInst_2_n3 ;
  wire   [63:0] StateRegOutput;
  wire   [31:0] AddConstOutput;
  wire   [47:0] Red_Plaintext;
  wire   [47:0] Red_StateRegOutput;
  wire   [23:0] Red_AddConstOutput;
  wire   [47:0] Red_ShiftRowsOutput;
  wire   [47:0] Red_Feedback;
  wire   [143:0] Red_SignaltoCheck;
  wire   [2:0] Error;
  wire   [3:0] \MCInst_MC0_v3_3 ;
  wire   [3:0] \MCInst_MC0_v3_2 ;
  wire   [3:0] \MCInst_MC0_v3_1 ;
  wire   [3:0] \MCInst_MC0_v3_0 ;
  wire   [3:0] \MCInst_MC0_v2_3 ;
  wire   [3:0] \MCInst_MC0_v2_2 ;
  wire   [3:0] \MCInst_MC0_v2_1 ;
  wire   [3:0] \MCInst_MC0_v2_0 ;
  wire   [3:0] \MCInst_MC0_v1_3 ;
  wire   [3:0] \MCInst_MC0_v1_2 ;
  wire   [3:0] \MCInst_MC0_v1_1 ;
  wire   [3:0] \MCInst_MC0_v1_0 ;
  wire   [3:0] \MCInst_MC0_v0_3 ;
  wire   [3:0] \MCInst_MC0_v0_2 ;
  wire   [3:0] \MCInst_MC0_v0_1 ;
  wire   [3:0] \MCInst_MC0_v0_0 ;
  wire   [3:0] \MCInst_MC1_v3_3 ;
  wire   [3:0] \MCInst_MC1_v3_2 ;
  wire   [3:0] \MCInst_MC1_v3_1 ;
  wire   [3:0] \MCInst_MC1_v3_0 ;
  wire   [3:0] \MCInst_MC1_v2_3 ;
  wire   [3:0] \MCInst_MC1_v2_2 ;
  wire   [3:0] \MCInst_MC1_v2_1 ;
  wire   [3:0] \MCInst_MC1_v2_0 ;
  wire   [3:0] \MCInst_MC1_v1_3 ;
  wire   [3:0] \MCInst_MC1_v1_2 ;
  wire   [3:0] \MCInst_MC1_v1_1 ;
  wire   [3:0] \MCInst_MC1_v1_0 ;
  wire   [3:0] \MCInst_MC1_v0_3 ;
  wire   [3:0] \MCInst_MC1_v0_2 ;
  wire   [3:0] \MCInst_MC1_v0_1 ;
  wire   [3:0] \MCInst_MC1_v0_0 ;
  wire   [3:0] \MCInst_MC2_v3_3 ;
  wire   [3:0] \MCInst_MC2_v3_2 ;
  wire   [3:0] \MCInst_MC2_v3_1 ;
  wire   [3:0] \MCInst_MC2_v3_0 ;
  wire   [3:0] \MCInst_MC2_v2_3 ;
  wire   [3:0] \MCInst_MC2_v2_2 ;
  wire   [3:0] \MCInst_MC2_v2_1 ;
  wire   [3:0] \MCInst_MC2_v2_0 ;
  wire   [3:0] \MCInst_MC2_v1_3 ;
  wire   [3:0] \MCInst_MC2_v1_2 ;
  wire   [3:0] \MCInst_MC2_v1_1 ;
  wire   [3:0] \MCInst_MC2_v1_0 ;
  wire   [3:0] \MCInst_MC2_v0_3 ;
  wire   [3:0] \MCInst_MC2_v0_2 ;
  wire   [3:0] \MCInst_MC2_v0_1 ;
  wire   [3:0] \MCInst_MC2_v0_0 ;
  wire   [3:0] \MCInst_MC3_v3_3 ;
  wire   [3:0] \MCInst_MC3_v3_2 ;
  wire   [3:0] \MCInst_MC3_v3_1 ;
  wire   [3:0] \MCInst_MC3_v3_0 ;
  wire   [3:0] \MCInst_MC3_v2_3 ;
  wire   [3:0] \MCInst_MC3_v2_2 ;
  wire   [3:0] \MCInst_MC3_v2_1 ;
  wire   [3:0] \MCInst_MC3_v2_0 ;
  wire   [3:0] \MCInst_MC3_v1_3 ;
  wire   [3:0] \MCInst_MC3_v1_2 ;
  wire   [3:0] \MCInst_MC3_v1_1 ;
  wire   [3:0] \MCInst_MC3_v1_0 ;
  wire   [3:0] \MCInst_MC3_v0_3 ;
  wire   [3:0] \MCInst_MC3_v0_2 ;
  wire   [3:0] \MCInst_MC3_v0_1 ;
  wire   [3:0] \MCInst_MC3_v0_0 ;
  wire   [2:0] \Red_MCInst_MC0_v3_3 ;
  wire   [2:0] \Red_MCInst_MC0_v3_2 ;
  wire   [2:0] \Red_MCInst_MC0_v3_1 ;
  wire   [2:0] \Red_MCInst_MC0_v3_0 ;
  wire   [2:0] \Red_MCInst_MC0_v2_3 ;
  wire   [2:0] \Red_MCInst_MC0_v2_2 ;
  wire   [2:0] \Red_MCInst_MC0_v2_1 ;
  wire   [2:0] \Red_MCInst_MC0_v2_0 ;
  wire   [2:0] \Red_MCInst_MC0_v1_3 ;
  wire   [2:0] \Red_MCInst_MC0_v1_2 ;
  wire   [2:0] \Red_MCInst_MC0_v1_1 ;
  wire   [2:0] \Red_MCInst_MC0_v1_0 ;
  wire   [2:0] \Red_MCInst_MC0_v0_3 ;
  wire   [2:0] \Red_MCInst_MC0_v0_2 ;
  wire   [2:0] \Red_MCInst_MC0_v0_1 ;
  wire   [2:0] \Red_MCInst_MC0_v0_0 ;
  wire   [2:0] \Red_MCInst_MC1_v3_3 ;
  wire   [2:0] \Red_MCInst_MC1_v3_2 ;
  wire   [2:0] \Red_MCInst_MC1_v3_1 ;
  wire   [2:0] \Red_MCInst_MC1_v3_0 ;
  wire   [2:0] \Red_MCInst_MC1_v2_3 ;
  wire   [2:0] \Red_MCInst_MC1_v2_2 ;
  wire   [2:0] \Red_MCInst_MC1_v2_1 ;
  wire   [2:0] \Red_MCInst_MC1_v2_0 ;
  wire   [2:0] \Red_MCInst_MC1_v1_3 ;
  wire   [2:0] \Red_MCInst_MC1_v1_2 ;
  wire   [2:0] \Red_MCInst_MC1_v1_1 ;
  wire   [2:0] \Red_MCInst_MC1_v1_0 ;
  wire   [2:0] \Red_MCInst_MC1_v0_3 ;
  wire   [2:0] \Red_MCInst_MC1_v0_2 ;
  wire   [2:0] \Red_MCInst_MC1_v0_1 ;
  wire   [2:0] \Red_MCInst_MC1_v0_0 ;
  wire   [2:0] \Red_MCInst_MC2_v3_3 ;
  wire   [2:0] \Red_MCInst_MC2_v3_2 ;
  wire   [2:0] \Red_MCInst_MC2_v3_1 ;
  wire   [2:0] \Red_MCInst_MC2_v3_0 ;
  wire   [2:0] \Red_MCInst_MC2_v2_3 ;
  wire   [2:0] \Red_MCInst_MC2_v2_2 ;
  wire   [2:0] \Red_MCInst_MC2_v2_1 ;
  wire   [2:0] \Red_MCInst_MC2_v2_0 ;
  wire   [2:0] \Red_MCInst_MC2_v1_3 ;
  wire   [2:0] \Red_MCInst_MC2_v1_2 ;
  wire   [2:0] \Red_MCInst_MC2_v1_1 ;
  wire   [2:0] \Red_MCInst_MC2_v1_0 ;
  wire   [2:0] \Red_MCInst_MC2_v0_3 ;
  wire   [2:0] \Red_MCInst_MC2_v0_2 ;
  wire   [2:0] \Red_MCInst_MC2_v0_1 ;
  wire   [2:0] \Red_MCInst_MC2_v0_0 ;
  wire   [2:0] \Red_MCInst_MC3_v3_3 ;
  wire   [2:0] \Red_MCInst_MC3_v3_2 ;
  wire   [2:0] \Red_MCInst_MC3_v3_1 ;
  wire   [2:0] \Red_MCInst_MC3_v3_0 ;
  wire   [2:0] \Red_MCInst_MC3_v2_3 ;
  wire   [2:0] \Red_MCInst_MC3_v2_2 ;
  wire   [2:0] \Red_MCInst_MC3_v2_1 ;
  wire   [2:0] \Red_MCInst_MC3_v2_0 ;
  wire   [2:0] \Red_MCInst_MC3_v1_3 ;
  wire   [2:0] \Red_MCInst_MC3_v1_2 ;
  wire   [2:0] \Red_MCInst_MC3_v1_1 ;
  wire   [2:0] \Red_MCInst_MC3_v1_0 ;
  wire   [2:0] \Red_MCInst_MC3_v0_3 ;
  wire   [2:0] \Red_MCInst_MC3_v0_2 ;
  wire   [2:0] \Red_MCInst_MC3_v0_1 ;
  wire   [2:0] \Red_MCInst_MC3_v0_0 ;

  AND2_X1 \Check1_CheckInst_U8 ( .A1(Error[2]), .A2(Error[0]), .ZN(n5) );
  NAND2_X1 \Check1_CheckInst_U9 ( .A1(Error[1]), .A2(n5), .ZN(ErrorFlag) );
  DFF_X1 \StateReg_s_current_state_reg[0]  ( .D(Plaintext[0]), .CK(clk), .Q(
        StateRegOutput[0]) );
  DFF_X1 \StateReg_s_current_state_reg[1]  ( .D(Plaintext[1]), .CK(clk), .Q(
        StateRegOutput[1]) );
  DFF_X1 \StateReg_s_current_state_reg[2]  ( .D(Plaintext[2]), .CK(clk), .Q(
        StateRegOutput[2]) );
  DFF_X1 \StateReg_s_current_state_reg[3]  ( .D(Plaintext[3]), .CK(clk), .Q(
        StateRegOutput[3]) );
  DFF_X1 \StateReg_s_current_state_reg[4]  ( .D(Plaintext[4]), .CK(clk), .Q(
        StateRegOutput[4]) );
  DFF_X1 \StateReg_s_current_state_reg[5]  ( .D(Plaintext[5]), .CK(clk), .Q(
        StateRegOutput[5]) );
  DFF_X1 \StateReg_s_current_state_reg[6]  ( .D(Plaintext[6]), .CK(clk), .Q(
        StateRegOutput[6]) );
  DFF_X1 \StateReg_s_current_state_reg[7]  ( .D(Plaintext[7]), .CK(clk), .Q(
        StateRegOutput[7]) );
  DFF_X1 \StateReg_s_current_state_reg[8]  ( .D(Plaintext[8]), .CK(clk), .Q(
        AddConstOutput[0]) );
  DFF_X1 \StateReg_s_current_state_reg[9]  ( .D(Plaintext[9]), .CK(clk), .Q(
        AddConstOutput[1]) );
  DFF_X1 \StateReg_s_current_state_reg[10]  ( .D(Plaintext[10]), .CK(clk), .Q(
        AddConstOutput[2]) );
  DFF_X1 \StateReg_s_current_state_reg[11]  ( .D(Plaintext[11]), .CK(clk), .Q(
        AddConstOutput[3]) );
  DFF_X1 \StateReg_s_current_state_reg[12]  ( .D(Plaintext[12]), .CK(clk), .Q(
        StateRegOutput[12]) );
  DFF_X1 \StateReg_s_current_state_reg[13]  ( .D(Plaintext[13]), .CK(clk), .Q(
        StateRegOutput[13]) );
  DFF_X1 \StateReg_s_current_state_reg[14]  ( .D(Plaintext[14]), .CK(clk), .Q(
        AddConstOutput[6]) );
  DFF_X1 \StateReg_s_current_state_reg[15]  ( .D(Plaintext[15]), .CK(clk), .Q(
        AddConstOutput[7]) );
  DFF_X1 \StateReg_s_current_state_reg[16]  ( .D(Plaintext[16]), .CK(clk), .Q(
        StateRegOutput[16]) );
  DFF_X1 \StateReg_s_current_state_reg[17]  ( .D(Plaintext[17]), .CK(clk), .Q(
        StateRegOutput[17]) );
  DFF_X1 \StateReg_s_current_state_reg[18]  ( .D(Plaintext[18]), .CK(clk), .Q(
        StateRegOutput[18]) );
  DFF_X1 \StateReg_s_current_state_reg[19]  ( .D(Plaintext[19]), .CK(clk), .Q(
        StateRegOutput[19]) );
  DFF_X1 \StateReg_s_current_state_reg[20]  ( .D(Plaintext[20]), .CK(clk), .Q(
        StateRegOutput[20]) );
  DFF_X1 \StateReg_s_current_state_reg[21]  ( .D(Plaintext[21]), .CK(clk), .Q(
        StateRegOutput[21]) );
  DFF_X1 \StateReg_s_current_state_reg[22]  ( .D(Plaintext[22]), .CK(clk), .Q(
        StateRegOutput[22]) );
  DFF_X1 \StateReg_s_current_state_reg[23]  ( .D(Plaintext[23]), .CK(clk), .Q(
        StateRegOutput[23]) );
  DFF_X1 \StateReg_s_current_state_reg[24]  ( .D(Plaintext[24]), .CK(clk), .Q(
        AddConstOutput[8]) );
  DFF_X1 \StateReg_s_current_state_reg[25]  ( .D(Plaintext[25]), .CK(clk), .Q(
        AddConstOutput[9]) );
  DFF_X1 \StateReg_s_current_state_reg[26]  ( .D(Plaintext[26]), .CK(clk), .Q(
        AddConstOutput[10]) );
  DFF_X1 \StateReg_s_current_state_reg[27]  ( .D(Plaintext[27]), .CK(clk), .Q(
        AddConstOutput[11]) );
  DFF_X1 \StateReg_s_current_state_reg[28]  ( .D(Plaintext[28]), .CK(clk), .Q(
        AddConstOutput[12]) );
  DFF_X1 \StateReg_s_current_state_reg[29]  ( .D(Plaintext[29]), .CK(clk), .Q(
        StateRegOutput[29]) );
  DFF_X1 \StateReg_s_current_state_reg[30]  ( .D(Plaintext[30]), .CK(clk), .Q(
        AddConstOutput[14]) );
  DFF_X1 \StateReg_s_current_state_reg[31]  ( .D(Plaintext[31]), .CK(clk), .Q(
        AddConstOutput[15]) );
  DFF_X1 \StateReg_s_current_state_reg[32]  ( .D(Plaintext[32]), .CK(clk), .Q(
        StateRegOutput[32]) );
  DFF_X1 \StateReg_s_current_state_reg[33]  ( .D(Plaintext[33]), .CK(clk), .Q(
        StateRegOutput[33]) );
  DFF_X1 \StateReg_s_current_state_reg[34]  ( .D(Plaintext[34]), .CK(clk), .Q(
        StateRegOutput[34]) );
  DFF_X1 \StateReg_s_current_state_reg[35]  ( .D(Plaintext[35]), .CK(clk), .Q(
        StateRegOutput[35]) );
  DFF_X1 \StateReg_s_current_state_reg[36]  ( .D(Plaintext[36]), .CK(clk), .Q(
        StateRegOutput[36]) );
  DFF_X1 \StateReg_s_current_state_reg[37]  ( .D(Plaintext[37]), .CK(clk), .Q(
        StateRegOutput[37]) );
  DFF_X1 \StateReg_s_current_state_reg[38]  ( .D(Plaintext[38]), .CK(clk), .Q(
        StateRegOutput[38]) );
  DFF_X1 \StateReg_s_current_state_reg[39]  ( .D(Plaintext[39]), .CK(clk), .Q(
        StateRegOutput[39]) );
  DFF_X1 \StateReg_s_current_state_reg[40]  ( .D(Plaintext[40]), .CK(clk), .Q(
        AddConstOutput[16]) );
  DFF_X1 \StateReg_s_current_state_reg[41]  ( .D(Plaintext[41]), .CK(clk), .Q(
        AddConstOutput[17]) );
  DFF_X1 \StateReg_s_current_state_reg[42]  ( .D(Plaintext[42]), .CK(clk), .Q(
        AddConstOutput[18]) );
  DFF_X1 \StateReg_s_current_state_reg[43]  ( .D(Plaintext[43]), .CK(clk), .Q(
        AddConstOutput[19]) );
  DFF_X1 \StateReg_s_current_state_reg[44]  ( .D(Plaintext[44]), .CK(clk), .Q(
        StateRegOutput[44]) );
  DFF_X1 \StateReg_s_current_state_reg[45]  ( .D(Plaintext[45]), .CK(clk), .Q(
        AddConstOutput[21]) );
  DFF_X1 \StateReg_s_current_state_reg[46]  ( .D(Plaintext[46]), .CK(clk), .Q(
        StateRegOutput[46]) );
  DFF_X1 \StateReg_s_current_state_reg[47]  ( .D(Plaintext[47]), .CK(clk), .Q(
        AddConstOutput[23]) );
  DFF_X1 \StateReg_s_current_state_reg[48]  ( .D(Plaintext[48]), .CK(clk), .Q(
        StateRegOutput[48]) );
  DFF_X1 \StateReg_s_current_state_reg[49]  ( .D(Plaintext[49]), .CK(clk), .Q(
        StateRegOutput[49]) );
  DFF_X1 \StateReg_s_current_state_reg[50]  ( .D(Plaintext[50]), .CK(clk), .Q(
        StateRegOutput[50]) );
  DFF_X1 \StateReg_s_current_state_reg[51]  ( .D(Plaintext[51]), .CK(clk), .Q(
        StateRegOutput[51]) );
  DFF_X1 \StateReg_s_current_state_reg[52]  ( .D(Plaintext[52]), .CK(clk), .Q(
        StateRegOutput[52]) );
  DFF_X1 \StateReg_s_current_state_reg[53]  ( .D(Plaintext[53]), .CK(clk), .Q(
        StateRegOutput[53]) );
  DFF_X1 \StateReg_s_current_state_reg[54]  ( .D(Plaintext[54]), .CK(clk), .Q(
        StateRegOutput[54]) );
  DFF_X1 \StateReg_s_current_state_reg[55]  ( .D(Plaintext[55]), .CK(clk), .Q(
        StateRegOutput[55]) );
  DFF_X1 \StateReg_s_current_state_reg[56]  ( .D(Plaintext[56]), .CK(clk), .Q(
        AddConstOutput[24]) );
  DFF_X1 \StateReg_s_current_state_reg[57]  ( .D(Plaintext[57]), .CK(clk), .Q(
        AddConstOutput[25]) );
  DFF_X1 \StateReg_s_current_state_reg[58]  ( .D(Plaintext[58]), .CK(clk), .Q(
        AddConstOutput[26]) );
  DFF_X1 \StateReg_s_current_state_reg[59]  ( .D(Plaintext[59]), .CK(clk), .Q(
        AddConstOutput[27]) );
  DFF_X1 \StateReg_s_current_state_reg[60]  ( .D(Plaintext[60]), .CK(clk), .Q(
        AddConstOutput[28]) );
  DFF_X1 \StateReg_s_current_state_reg[61]  ( .D(Plaintext[61]), .CK(clk), .Q(
        AddConstOutput[29]) );
  DFF_X1 \StateReg_s_current_state_reg[62]  ( .D(Plaintext[62]), .CK(clk), .Q(
        StateRegOutput[62]) );
  DFF_X1 \StateReg_s_current_state_reg[63]  ( .D(Plaintext[63]), .CK(clk), .Q(
        AddConstOutput[31]) );
  INV_X1 \AddConstXOR_XORInst_XORInst_1_0_U1  ( .A(StateRegOutput[12]), .ZN(
        AddConstOutput[4]) );
  INV_X1 \AddConstXOR_XORInst_XORInst_1_1_U1  ( .A(StateRegOutput[13]), .ZN(
        AddConstOutput[5]) );
  INV_X1 \AddConstXOR_XORInst_XORInst_3_1_U1  ( .A(StateRegOutput[29]), .ZN(
        AddConstOutput[13]) );
  INV_X1 \AddConstXOR_XORInst_XORInst_5_0_U1  ( .A(StateRegOutput[44]), .ZN(
        AddConstOutput[20]) );
  INV_X1 \AddConstXOR_XORInst_XORInst_5_2_U1  ( .A(StateRegOutput[46]), .ZN(
        AddConstOutput[22]) );
  INV_X1 \AddConstXOR_XORInst_XORInst_7_2_U1  ( .A(StateRegOutput[62]), .ZN(
        AddConstOutput[30]) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_0_U7  ( .A1(StateRegOutput[2]), .A2(
        \SubCellInst_LFInst_0_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_0_LFInst_0_U6  ( .A(StateRegOutput[1]), .ZN(
        \SubCellInst_LFInst_0_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_0_LFInst_0_U5  ( .A(StateRegOutput[0]), .B(
        StateRegOutput[3]), .Z(\SubCellInst_LFInst_0_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_0_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_0_LFInst_0_n10 ), .ZN(\MCInst_MC0_v3_2 [3]) );
  XOR2_X1 \SubCellInst_LFInst_0_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_0_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_0_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_0_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_0_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_0_LFInst_1_n17 ), .ZN(\Red_MCInst_MC0_v3_3 [2]) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U11  ( .A1(StateRegOutput[1]), .A2(
        \SubCellInst_LFInst_0_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_1_U10  ( .A1(StateRegOutput[3]), .A2(
        \SubCellInst_LFInst_0_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_0_LFInst_1_U9  ( .A1(StateRegOutput[0]), .A2(
        StateRegOutput[2]), .ZN(\SubCellInst_LFInst_0_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U8  ( .A1(StateRegOutput[3]), .A2(
        \SubCellInst_LFInst_0_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_0_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_0_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U6  ( .A1(StateRegOutput[0]), .A2(
        StateRegOutput[2]), .ZN(\SubCellInst_LFInst_0_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_0_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_0_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U4  ( .A1(StateRegOutput[0]), .A2(
        StateRegOutput[1]), .ZN(\SubCellInst_LFInst_0_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_0_LFInst_1_U3  ( .A(StateRegOutput[2]), .ZN(
        \SubCellInst_LFInst_0_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_0_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_0_LFInst_2_n21 ), .ZN(\MCInst_MC0_v3_0 [3]) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U10  ( .A1(StateRegOutput[2]), .A2(
        \SubCellInst_LFInst_0_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_2_U9  ( .A1(StateRegOutput[1]), .A2(
        \SubCellInst_LFInst_0_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_0_LFInst_2_U8  ( .A(StateRegOutput[3]), .ZN(
        \SubCellInst_LFInst_0_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_0_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_0_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_0_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_0_LFInst_2_n16 ), .B(StateRegOutput[2]), .Z(
        \SubCellInst_LFInst_0_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U5  ( .A1(StateRegOutput[0]), .A2(
        StateRegOutput[1]), .ZN(\SubCellInst_LFInst_0_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_0_LFInst_2_n15 ), .A2(StateRegOutput[3]), .ZN(
        \SubCellInst_LFInst_0_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_0_LFInst_2_U3  ( .A(StateRegOutput[0]), .B(
        StateRegOutput[1]), .ZN(\SubCellInst_LFInst_0_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_0_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_0_LFInst_3_n15 ), .ZN(\Red_MCInst_MC0_v3_1 [2]) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_3_U8  ( .A1(StateRegOutput[1]), .A2(
        \SubCellInst_LFInst_0_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_0_LFInst_3_U7  ( .A(StateRegOutput[3]), .B(
        StateRegOutput[2]), .Z(\SubCellInst_LFInst_0_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_0_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_0_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_3_U5  ( .A1(StateRegOutput[0]), .A2(
        StateRegOutput[2]), .ZN(\SubCellInst_LFInst_0_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_0_LFInst_3_U4  ( .A(StateRegOutput[0]), .B(
        \SubCellInst_LFInst_0_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_0_LFInst_3_U3  ( .A1(StateRegOutput[3]), .A2(
        StateRegOutput[1]), .ZN(\SubCellInst_LFInst_0_LFInst_3_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_0_U7  ( .A1(StateRegOutput[6]), .A2(
        \SubCellInst_LFInst_1_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_1_LFInst_0_U6  ( .A(StateRegOutput[5]), .ZN(
        \SubCellInst_LFInst_1_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_1_LFInst_0_U5  ( .A(StateRegOutput[4]), .B(
        StateRegOutput[7]), .Z(\SubCellInst_LFInst_1_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_1_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_1_LFInst_0_n10 ), .ZN(\MCInst_MC3_v3_2 [3]) );
  XOR2_X1 \SubCellInst_LFInst_1_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_1_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_1_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_1_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_1_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_1_LFInst_1_n17 ), .ZN(\Red_MCInst_MC3_v3_3 [2]) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U11  ( .A1(StateRegOutput[5]), .A2(
        \SubCellInst_LFInst_1_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_1_U10  ( .A1(StateRegOutput[7]), .A2(
        \SubCellInst_LFInst_1_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_1_LFInst_1_U9  ( .A1(StateRegOutput[4]), .A2(
        StateRegOutput[6]), .ZN(\SubCellInst_LFInst_1_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U8  ( .A1(StateRegOutput[7]), .A2(
        \SubCellInst_LFInst_1_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_1_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_1_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U6  ( .A1(StateRegOutput[4]), .A2(
        StateRegOutput[6]), .ZN(\SubCellInst_LFInst_1_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_1_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_1_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U4  ( .A1(StateRegOutput[4]), .A2(
        StateRegOutput[5]), .ZN(\SubCellInst_LFInst_1_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_1_LFInst_1_U3  ( .A(StateRegOutput[6]), .ZN(
        \SubCellInst_LFInst_1_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_1_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_1_LFInst_2_n21 ), .ZN(\MCInst_MC3_v3_0 [3]) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U10  ( .A1(StateRegOutput[6]), .A2(
        \SubCellInst_LFInst_1_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_2_U9  ( .A1(StateRegOutput[5]), .A2(
        \SubCellInst_LFInst_1_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_1_LFInst_2_U8  ( .A(StateRegOutput[7]), .ZN(
        \SubCellInst_LFInst_1_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_1_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_1_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_1_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_1_LFInst_2_n16 ), .B(StateRegOutput[6]), .Z(
        \SubCellInst_LFInst_1_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U5  ( .A1(StateRegOutput[4]), .A2(
        StateRegOutput[5]), .ZN(\SubCellInst_LFInst_1_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_1_LFInst_2_n15 ), .A2(StateRegOutput[7]), .ZN(
        \SubCellInst_LFInst_1_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_1_LFInst_2_U3  ( .A(StateRegOutput[4]), .B(
        StateRegOutput[5]), .ZN(\SubCellInst_LFInst_1_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_1_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_1_LFInst_3_n15 ), .ZN(\Red_MCInst_MC3_v3_1 [2]) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_3_U8  ( .A1(StateRegOutput[5]), .A2(
        \SubCellInst_LFInst_1_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_1_LFInst_3_U7  ( .A(StateRegOutput[7]), .B(
        StateRegOutput[6]), .Z(\SubCellInst_LFInst_1_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_1_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_1_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_3_U5  ( .A1(StateRegOutput[4]), .A2(
        StateRegOutput[6]), .ZN(\SubCellInst_LFInst_1_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_1_LFInst_3_U4  ( .A(StateRegOutput[4]), .B(
        \SubCellInst_LFInst_1_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_1_LFInst_3_U3  ( .A1(StateRegOutput[7]), .A2(
        StateRegOutput[5]), .ZN(\SubCellInst_LFInst_1_LFInst_3_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_0_U7  ( .A1(AddConstOutput[2]), .A2(
        \SubCellInst_LFInst_2_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_2_LFInst_0_U6  ( .A(AddConstOutput[1]), .ZN(
        \SubCellInst_LFInst_2_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_2_LFInst_0_U5  ( .A(AddConstOutput[0]), .B(
        AddConstOutput[3]), .Z(\SubCellInst_LFInst_2_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_2_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_2_LFInst_0_n10 ), .ZN(\MCInst_MC2_v3_2 [3]) );
  XOR2_X1 \SubCellInst_LFInst_2_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_2_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_2_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_2_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_2_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_2_LFInst_1_n17 ), .ZN(\Red_MCInst_MC2_v3_3 [2]) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U11  ( .A1(AddConstOutput[1]), .A2(
        \SubCellInst_LFInst_2_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_1_U10  ( .A1(AddConstOutput[3]), .A2(
        \SubCellInst_LFInst_2_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_2_LFInst_1_U9  ( .A1(AddConstOutput[0]), .A2(
        AddConstOutput[2]), .ZN(\SubCellInst_LFInst_2_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U8  ( .A1(AddConstOutput[3]), .A2(
        \SubCellInst_LFInst_2_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_2_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_2_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U6  ( .A1(AddConstOutput[0]), .A2(
        AddConstOutput[2]), .ZN(\SubCellInst_LFInst_2_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_2_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_2_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U4  ( .A1(AddConstOutput[0]), .A2(
        AddConstOutput[1]), .ZN(\SubCellInst_LFInst_2_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_2_LFInst_1_U3  ( .A(AddConstOutput[2]), .ZN(
        \SubCellInst_LFInst_2_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_2_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_2_LFInst_2_n21 ), .ZN(\MCInst_MC2_v3_0 [3]) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U10  ( .A1(AddConstOutput[2]), .A2(
        \SubCellInst_LFInst_2_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_2_U9  ( .A1(AddConstOutput[1]), .A2(
        \SubCellInst_LFInst_2_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_2_LFInst_2_U8  ( .A(AddConstOutput[3]), .ZN(
        \SubCellInst_LFInst_2_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_2_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_2_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_2_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_2_LFInst_2_n16 ), .B(AddConstOutput[2]), .Z(
        \SubCellInst_LFInst_2_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U5  ( .A1(AddConstOutput[0]), .A2(
        AddConstOutput[1]), .ZN(\SubCellInst_LFInst_2_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_2_LFInst_2_n15 ), .A2(AddConstOutput[3]), .ZN(
        \SubCellInst_LFInst_2_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_2_LFInst_2_U3  ( .A(AddConstOutput[0]), .B(
        AddConstOutput[1]), .ZN(\SubCellInst_LFInst_2_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_2_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_2_LFInst_3_n15 ), .ZN(\Red_MCInst_MC2_v3_1 [2]) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_3_U8  ( .A1(AddConstOutput[1]), .A2(
        \SubCellInst_LFInst_2_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_2_LFInst_3_U7  ( .A(AddConstOutput[3]), .B(
        AddConstOutput[2]), .Z(\SubCellInst_LFInst_2_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_2_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_2_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_3_U5  ( .A1(AddConstOutput[0]), .A2(
        AddConstOutput[2]), .ZN(\SubCellInst_LFInst_2_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_2_LFInst_3_U4  ( .A(AddConstOutput[0]), .B(
        \SubCellInst_LFInst_2_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_2_LFInst_3_U3  ( .A1(AddConstOutput[3]), .A2(
        AddConstOutput[1]), .ZN(\SubCellInst_LFInst_2_LFInst_3_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_0_U7  ( .A1(AddConstOutput[6]), .A2(
        \SubCellInst_LFInst_3_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_3_LFInst_0_U6  ( .A(AddConstOutput[5]), .ZN(
        \SubCellInst_LFInst_3_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_3_LFInst_0_U5  ( .A(AddConstOutput[4]), .B(
        AddConstOutput[7]), .Z(\SubCellInst_LFInst_3_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_3_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_3_LFInst_0_n10 ), .ZN(\MCInst_MC1_v3_2 [3]) );
  XOR2_X1 \SubCellInst_LFInst_3_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_3_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_3_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_3_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_3_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_3_LFInst_1_n17 ), .ZN(\Red_MCInst_MC1_v3_3 [2]) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U11  ( .A1(AddConstOutput[5]), .A2(
        \SubCellInst_LFInst_3_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_1_U10  ( .A1(AddConstOutput[7]), .A2(
        \SubCellInst_LFInst_3_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_3_LFInst_1_U9  ( .A1(AddConstOutput[4]), .A2(
        AddConstOutput[6]), .ZN(\SubCellInst_LFInst_3_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U8  ( .A1(AddConstOutput[7]), .A2(
        \SubCellInst_LFInst_3_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_3_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_3_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U6  ( .A1(AddConstOutput[4]), .A2(
        AddConstOutput[6]), .ZN(\SubCellInst_LFInst_3_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_3_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_3_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U4  ( .A1(AddConstOutput[4]), .A2(
        AddConstOutput[5]), .ZN(\SubCellInst_LFInst_3_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_3_LFInst_1_U3  ( .A(AddConstOutput[6]), .ZN(
        \SubCellInst_LFInst_3_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_3_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_3_LFInst_2_n21 ), .ZN(\MCInst_MC1_v3_0 [3]) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U10  ( .A1(AddConstOutput[6]), .A2(
        \SubCellInst_LFInst_3_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_2_U9  ( .A1(AddConstOutput[5]), .A2(
        \SubCellInst_LFInst_3_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_3_LFInst_2_U8  ( .A(AddConstOutput[7]), .ZN(
        \SubCellInst_LFInst_3_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_3_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_3_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_3_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_3_LFInst_2_n16 ), .B(AddConstOutput[6]), .Z(
        \SubCellInst_LFInst_3_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U5  ( .A1(AddConstOutput[4]), .A2(
        AddConstOutput[5]), .ZN(\SubCellInst_LFInst_3_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_3_LFInst_2_n15 ), .A2(AddConstOutput[7]), .ZN(
        \SubCellInst_LFInst_3_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_3_LFInst_2_U3  ( .A(AddConstOutput[4]), .B(
        AddConstOutput[5]), .ZN(\SubCellInst_LFInst_3_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_3_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_3_LFInst_3_n15 ), .ZN(\Red_MCInst_MC1_v3_1 [2]) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_3_U8  ( .A1(AddConstOutput[5]), .A2(
        \SubCellInst_LFInst_3_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_3_LFInst_3_U7  ( .A(AddConstOutput[7]), .B(
        AddConstOutput[6]), .Z(\SubCellInst_LFInst_3_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_3_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_3_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_3_U5  ( .A1(AddConstOutput[4]), .A2(
        AddConstOutput[6]), .ZN(\SubCellInst_LFInst_3_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_3_LFInst_3_U4  ( .A(AddConstOutput[4]), .B(
        \SubCellInst_LFInst_3_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_3_LFInst_3_U3  ( .A1(AddConstOutput[7]), .A2(
        AddConstOutput[5]), .ZN(\SubCellInst_LFInst_3_LFInst_3_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_0_U7  ( .A1(StateRegOutput[18]), .A2(
        \SubCellInst_LFInst_4_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_4_LFInst_0_U6  ( .A(StateRegOutput[17]), .ZN(
        \SubCellInst_LFInst_4_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_4_LFInst_0_U5  ( .A(StateRegOutput[16]), .B(
        StateRegOutput[19]), .Z(\SubCellInst_LFInst_4_LFInst_0_n9 ) );
  INV_X2 \SubCellInst_LFInst_4_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_4_LFInst_0_n10 ), .ZN(\Red_MCInst_MC1_v2_1 [1]) );
  XOR2_X1 \SubCellInst_LFInst_4_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_4_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_4_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_4_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_4_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_4_LFInst_1_n17 ), .ZN(\MCInst_MC1_v2_0 [2]) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U11  ( .A1(StateRegOutput[17]), .A2(
        \SubCellInst_LFInst_4_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_1_U10  ( .A1(StateRegOutput[19]), .A2(
        \SubCellInst_LFInst_4_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_4_LFInst_1_U9  ( .A1(StateRegOutput[16]), .A2(
        StateRegOutput[18]), .ZN(\SubCellInst_LFInst_4_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U8  ( .A1(StateRegOutput[19]), .A2(
        \SubCellInst_LFInst_4_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_4_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_4_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U6  ( .A1(StateRegOutput[16]), .A2(
        StateRegOutput[18]), .ZN(\SubCellInst_LFInst_4_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_4_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_4_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U4  ( .A1(StateRegOutput[16]), .A2(
        StateRegOutput[17]), .ZN(\SubCellInst_LFInst_4_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_4_LFInst_1_U3  ( .A(StateRegOutput[18]), .ZN(
        \SubCellInst_LFInst_4_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_4_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_4_LFInst_2_n21 ), .ZN(\MCInst_MC1_v2_0 [3]) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U10  ( .A1(StateRegOutput[18]), .A2(
        \SubCellInst_LFInst_4_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_2_U9  ( .A1(StateRegOutput[17]), .A2(
        \SubCellInst_LFInst_4_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_4_LFInst_2_U8  ( .A(StateRegOutput[19]), .ZN(
        \SubCellInst_LFInst_4_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_4_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_4_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_4_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_4_LFInst_2_n16 ), .B(StateRegOutput[18]), .Z(
        \SubCellInst_LFInst_4_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U5  ( .A1(StateRegOutput[16]), .A2(
        StateRegOutput[17]), .ZN(\SubCellInst_LFInst_4_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_4_LFInst_2_n15 ), .A2(StateRegOutput[19]), .ZN(
        \SubCellInst_LFInst_4_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_4_LFInst_2_U3  ( .A(StateRegOutput[16]), .B(
        StateRegOutput[17]), .ZN(\SubCellInst_LFInst_4_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_3_U9  ( .A1(StateRegOutput[17]), .A2(
        \SubCellInst_LFInst_4_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_4_LFInst_3_U8  ( .A(StateRegOutput[19]), .B(
        StateRegOutput[18]), .Z(\SubCellInst_LFInst_4_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_3_U7  ( .A1(
        \SubCellInst_LFInst_4_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_4_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_3_U6  ( .A1(StateRegOutput[16]), .A2(
        StateRegOutput[18]), .ZN(\SubCellInst_LFInst_4_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_4_LFInst_3_U5  ( .A(StateRegOutput[16]), .B(
        \SubCellInst_LFInst_4_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_4_LFInst_3_U4  ( .A1(StateRegOutput[19]), .A2(
        StateRegOutput[17]), .ZN(\SubCellInst_LFInst_4_LFInst_3_n11 ) );
  NAND2_X2 \SubCellInst_LFInst_4_LFInst_3_U3  ( .A1(
        \SubCellInst_LFInst_4_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_4_LFInst_3_n15 ), .ZN(\Red_MCInst_MC1_v2_2 [1]) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_0_U7  ( .A1(StateRegOutput[22]), .A2(
        \SubCellInst_LFInst_5_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_5_LFInst_0_U6  ( .A(StateRegOutput[21]), .ZN(
        \SubCellInst_LFInst_5_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_5_LFInst_0_U5  ( .A(StateRegOutput[20]), .B(
        StateRegOutput[23]), .Z(\SubCellInst_LFInst_5_LFInst_0_n9 ) );
  INV_X2 \SubCellInst_LFInst_5_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_5_LFInst_0_n10 ), .ZN(\Red_MCInst_MC0_v2_1 [1]) );
  XOR2_X1 \SubCellInst_LFInst_5_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_5_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_5_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_5_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_5_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_5_LFInst_1_n17 ), .ZN(\MCInst_MC0_v2_0 [2]) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U11  ( .A1(StateRegOutput[21]), .A2(
        \SubCellInst_LFInst_5_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_1_U10  ( .A1(StateRegOutput[23]), .A2(
        \SubCellInst_LFInst_5_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_5_LFInst_1_U9  ( .A1(StateRegOutput[20]), .A2(
        StateRegOutput[22]), .ZN(\SubCellInst_LFInst_5_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U8  ( .A1(StateRegOutput[23]), .A2(
        \SubCellInst_LFInst_5_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_5_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_5_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U6  ( .A1(StateRegOutput[20]), .A2(
        StateRegOutput[22]), .ZN(\SubCellInst_LFInst_5_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_5_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_5_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U4  ( .A1(StateRegOutput[20]), .A2(
        StateRegOutput[21]), .ZN(\SubCellInst_LFInst_5_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_5_LFInst_1_U3  ( .A(StateRegOutput[22]), .ZN(
        \SubCellInst_LFInst_5_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_5_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_5_LFInst_2_n21 ), .ZN(\MCInst_MC0_v2_0 [3]) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U10  ( .A1(StateRegOutput[22]), .A2(
        \SubCellInst_LFInst_5_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_2_U9  ( .A1(StateRegOutput[21]), .A2(
        \SubCellInst_LFInst_5_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_5_LFInst_2_U8  ( .A(StateRegOutput[23]), .ZN(
        \SubCellInst_LFInst_5_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_5_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_5_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_5_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_5_LFInst_2_n16 ), .B(StateRegOutput[22]), .Z(
        \SubCellInst_LFInst_5_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U5  ( .A1(StateRegOutput[20]), .A2(
        StateRegOutput[21]), .ZN(\SubCellInst_LFInst_5_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_5_LFInst_2_n15 ), .A2(StateRegOutput[23]), .ZN(
        \SubCellInst_LFInst_5_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_5_LFInst_2_U3  ( .A(StateRegOutput[20]), .B(
        StateRegOutput[21]), .ZN(\SubCellInst_LFInst_5_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_3_U9  ( .A1(StateRegOutput[21]), .A2(
        \SubCellInst_LFInst_5_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_5_LFInst_3_U8  ( .A(StateRegOutput[23]), .B(
        StateRegOutput[22]), .Z(\SubCellInst_LFInst_5_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_3_U7  ( .A1(
        \SubCellInst_LFInst_5_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_5_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_3_U6  ( .A1(StateRegOutput[20]), .A2(
        StateRegOutput[22]), .ZN(\SubCellInst_LFInst_5_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_5_LFInst_3_U5  ( .A(StateRegOutput[20]), .B(
        \SubCellInst_LFInst_5_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_5_LFInst_3_U4  ( .A1(StateRegOutput[23]), .A2(
        StateRegOutput[21]), .ZN(\SubCellInst_LFInst_5_LFInst_3_n11 ) );
  NAND2_X2 \SubCellInst_LFInst_5_LFInst_3_U3  ( .A1(
        \SubCellInst_LFInst_5_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_5_LFInst_3_n15 ), .ZN(\Red_MCInst_MC0_v2_2 [1]) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_0_U7  ( .A1(AddConstOutput[10]), .A2(
        \SubCellInst_LFInst_6_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_6_LFInst_0_U6  ( .A(AddConstOutput[9]), .ZN(
        \SubCellInst_LFInst_6_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_6_LFInst_0_U5  ( .A(AddConstOutput[8]), .B(
        AddConstOutput[11]), .Z(\SubCellInst_LFInst_6_LFInst_0_n9 ) );
  INV_X2 \SubCellInst_LFInst_6_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_6_LFInst_0_n10 ), .ZN(\Red_MCInst_MC3_v2_1 [1]) );
  XOR2_X1 \SubCellInst_LFInst_6_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_6_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_6_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_6_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_6_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_6_LFInst_1_n17 ), .ZN(\MCInst_MC3_v2_0 [2]) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U11  ( .A1(AddConstOutput[9]), .A2(
        \SubCellInst_LFInst_6_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_1_U10  ( .A1(AddConstOutput[11]), .A2(
        \SubCellInst_LFInst_6_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_6_LFInst_1_U9  ( .A1(AddConstOutput[8]), .A2(
        AddConstOutput[10]), .ZN(\SubCellInst_LFInst_6_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U8  ( .A1(AddConstOutput[11]), .A2(
        \SubCellInst_LFInst_6_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_6_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_6_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U6  ( .A1(AddConstOutput[8]), .A2(
        AddConstOutput[10]), .ZN(\SubCellInst_LFInst_6_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_6_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_6_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U4  ( .A1(AddConstOutput[8]), .A2(
        AddConstOutput[9]), .ZN(\SubCellInst_LFInst_6_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_6_LFInst_1_U3  ( .A(AddConstOutput[10]), .ZN(
        \SubCellInst_LFInst_6_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_6_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_6_LFInst_2_n21 ), .ZN(\MCInst_MC3_v2_0 [3]) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U10  ( .A1(AddConstOutput[10]), .A2(
        \SubCellInst_LFInst_6_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_2_U9  ( .A1(AddConstOutput[9]), .A2(
        \SubCellInst_LFInst_6_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_6_LFInst_2_U8  ( .A(AddConstOutput[11]), .ZN(
        \SubCellInst_LFInst_6_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_6_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_6_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_6_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_6_LFInst_2_n16 ), .B(AddConstOutput[10]), .Z(
        \SubCellInst_LFInst_6_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U5  ( .A1(AddConstOutput[8]), .A2(
        AddConstOutput[9]), .ZN(\SubCellInst_LFInst_6_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_6_LFInst_2_n15 ), .A2(AddConstOutput[11]), .ZN(
        \SubCellInst_LFInst_6_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_6_LFInst_2_U3  ( .A(AddConstOutput[8]), .B(
        AddConstOutput[9]), .ZN(\SubCellInst_LFInst_6_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_3_U9  ( .A1(AddConstOutput[9]), .A2(
        \SubCellInst_LFInst_6_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_6_LFInst_3_U8  ( .A(AddConstOutput[11]), .B(
        AddConstOutput[10]), .Z(\SubCellInst_LFInst_6_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_3_U7  ( .A1(
        \SubCellInst_LFInst_6_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_6_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_3_U6  ( .A1(AddConstOutput[8]), .A2(
        AddConstOutput[10]), .ZN(\SubCellInst_LFInst_6_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_6_LFInst_3_U5  ( .A(AddConstOutput[8]), .B(
        \SubCellInst_LFInst_6_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_6_LFInst_3_U4  ( .A1(AddConstOutput[11]), .A2(
        AddConstOutput[9]), .ZN(\SubCellInst_LFInst_6_LFInst_3_n11 ) );
  NAND2_X2 \SubCellInst_LFInst_6_LFInst_3_U3  ( .A1(
        \SubCellInst_LFInst_6_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_6_LFInst_3_n15 ), .ZN(\Red_MCInst_MC3_v2_2 [1]) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_0_U7  ( .A1(AddConstOutput[14]), .A2(
        \SubCellInst_LFInst_7_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_7_LFInst_0_U6  ( .A(AddConstOutput[13]), .ZN(
        \SubCellInst_LFInst_7_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_7_LFInst_0_U5  ( .A(AddConstOutput[12]), .B(
        AddConstOutput[15]), .Z(\SubCellInst_LFInst_7_LFInst_0_n9 ) );
  INV_X2 \SubCellInst_LFInst_7_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_7_LFInst_0_n10 ), .ZN(\Red_MCInst_MC2_v2_1 [1]) );
  XOR2_X1 \SubCellInst_LFInst_7_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_7_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_7_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_7_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_7_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_7_LFInst_1_n17 ), .ZN(\MCInst_MC2_v2_0 [2]) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U11  ( .A1(AddConstOutput[13]), .A2(
        \SubCellInst_LFInst_7_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_1_U10  ( .A1(AddConstOutput[15]), .A2(
        \SubCellInst_LFInst_7_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_7_LFInst_1_U9  ( .A1(AddConstOutput[12]), .A2(
        AddConstOutput[14]), .ZN(\SubCellInst_LFInst_7_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U8  ( .A1(AddConstOutput[15]), .A2(
        \SubCellInst_LFInst_7_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_7_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_7_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U6  ( .A1(AddConstOutput[12]), .A2(
        AddConstOutput[14]), .ZN(\SubCellInst_LFInst_7_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_7_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_7_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U4  ( .A1(AddConstOutput[12]), .A2(
        AddConstOutput[13]), .ZN(\SubCellInst_LFInst_7_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_7_LFInst_1_U3  ( .A(AddConstOutput[14]), .ZN(
        \SubCellInst_LFInst_7_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_7_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_7_LFInst_2_n21 ), .ZN(\MCInst_MC2_v2_0 [3]) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U10  ( .A1(AddConstOutput[14]), .A2(
        \SubCellInst_LFInst_7_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_2_U9  ( .A1(AddConstOutput[13]), .A2(
        \SubCellInst_LFInst_7_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_7_LFInst_2_U8  ( .A(AddConstOutput[15]), .ZN(
        \SubCellInst_LFInst_7_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_7_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_7_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_7_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_7_LFInst_2_n16 ), .B(AddConstOutput[14]), .Z(
        \SubCellInst_LFInst_7_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U5  ( .A1(AddConstOutput[12]), .A2(
        AddConstOutput[13]), .ZN(\SubCellInst_LFInst_7_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_7_LFInst_2_n15 ), .A2(AddConstOutput[15]), .ZN(
        \SubCellInst_LFInst_7_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_7_LFInst_2_U3  ( .A(AddConstOutput[12]), .B(
        AddConstOutput[13]), .ZN(\SubCellInst_LFInst_7_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_3_U9  ( .A1(AddConstOutput[13]), .A2(
        \SubCellInst_LFInst_7_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_7_LFInst_3_U8  ( .A(AddConstOutput[15]), .B(
        AddConstOutput[14]), .Z(\SubCellInst_LFInst_7_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_3_U7  ( .A1(
        \SubCellInst_LFInst_7_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_7_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_3_U6  ( .A1(AddConstOutput[12]), .A2(
        AddConstOutput[14]), .ZN(\SubCellInst_LFInst_7_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_7_LFInst_3_U5  ( .A(AddConstOutput[12]), .B(
        \SubCellInst_LFInst_7_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_7_LFInst_3_U4  ( .A1(AddConstOutput[15]), .A2(
        AddConstOutput[13]), .ZN(\SubCellInst_LFInst_7_LFInst_3_n11 ) );
  NAND2_X2 \SubCellInst_LFInst_7_LFInst_3_U3  ( .A1(
        \SubCellInst_LFInst_7_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_7_LFInst_3_n15 ), .ZN(\Red_MCInst_MC2_v2_2 [1]) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_0_U7  ( .A1(StateRegOutput[34]), .A2(
        \SubCellInst_LFInst_8_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_8_LFInst_0_U6  ( .A(StateRegOutput[33]), .ZN(
        \SubCellInst_LFInst_8_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_8_LFInst_0_U5  ( .A(StateRegOutput[32]), .B(
        StateRegOutput[35]), .Z(\SubCellInst_LFInst_8_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_8_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_8_LFInst_0_n10 ), .ZN(\MCInst_MC2_v1_0 [0]) );
  XOR2_X1 \SubCellInst_LFInst_8_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_8_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_8_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_8_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_1_U12  ( .A1(StateRegOutput[33]), .A2(
        \SubCellInst_LFInst_8_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_1_U11  ( .A1(StateRegOutput[35]), .A2(
        \SubCellInst_LFInst_8_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_8_LFInst_1_U10  ( .A1(StateRegOutput[32]), .A2(
        StateRegOutput[34]), .ZN(\SubCellInst_LFInst_8_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_1_U9  ( .A1(StateRegOutput[35]), .A2(
        \SubCellInst_LFInst_8_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_1_U8  ( .A1(
        \SubCellInst_LFInst_8_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_8_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_1_U7  ( .A1(StateRegOutput[32]), .A2(
        StateRegOutput[34]), .ZN(\SubCellInst_LFInst_8_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_8_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_8_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_1_U5  ( .A1(StateRegOutput[32]), .A2(
        StateRegOutput[33]), .ZN(\SubCellInst_LFInst_8_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_8_LFInst_1_U4  ( .A(StateRegOutput[34]), .ZN(
        \SubCellInst_LFInst_8_LFInst_1_n11 ) );
  NAND2_X2 \SubCellInst_LFInst_8_LFInst_1_U3  ( .A1(
        \SubCellInst_LFInst_8_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_8_LFInst_1_n17 ), .ZN(\Red_MCInst_MC2_v1_2 [1]) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_8_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_8_LFInst_2_n21 ), .ZN(\MCInst_MC2_v1_3 [3]) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U10  ( .A1(StateRegOutput[34]), .A2(
        \SubCellInst_LFInst_8_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_2_U9  ( .A1(StateRegOutput[33]), .A2(
        \SubCellInst_LFInst_8_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_8_LFInst_2_U8  ( .A(StateRegOutput[35]), .ZN(
        \SubCellInst_LFInst_8_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_8_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_8_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_8_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_8_LFInst_2_n16 ), .B(StateRegOutput[34]), .Z(
        \SubCellInst_LFInst_8_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U5  ( .A1(StateRegOutput[32]), .A2(
        StateRegOutput[33]), .ZN(\SubCellInst_LFInst_8_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_8_LFInst_2_n15 ), .A2(StateRegOutput[35]), .ZN(
        \SubCellInst_LFInst_8_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_8_LFInst_2_U3  ( .A(StateRegOutput[32]), .B(
        StateRegOutput[33]), .ZN(\SubCellInst_LFInst_8_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_8_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_8_LFInst_3_n15 ), .ZN(\Red_MCInst_MC2_v1_1 [2]) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_3_U8  ( .A1(StateRegOutput[33]), .A2(
        \SubCellInst_LFInst_8_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_8_LFInst_3_U7  ( .A(StateRegOutput[35]), .B(
        StateRegOutput[34]), .Z(\SubCellInst_LFInst_8_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_8_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_8_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_3_U5  ( .A1(StateRegOutput[32]), .A2(
        StateRegOutput[34]), .ZN(\SubCellInst_LFInst_8_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_8_LFInst_3_U4  ( .A(StateRegOutput[32]), .B(
        \SubCellInst_LFInst_8_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_8_LFInst_3_U3  ( .A1(StateRegOutput[35]), .A2(
        StateRegOutput[33]), .ZN(\SubCellInst_LFInst_8_LFInst_3_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_0_U7  ( .A1(StateRegOutput[38]), .A2(
        \SubCellInst_LFInst_9_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_9_LFInst_0_U6  ( .A(StateRegOutput[37]), .ZN(
        \SubCellInst_LFInst_9_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_9_LFInst_0_U5  ( .A(StateRegOutput[36]), .B(
        StateRegOutput[39]), .Z(\SubCellInst_LFInst_9_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_9_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_9_LFInst_0_n10 ), .ZN(\MCInst_MC1_v1_0 [0]) );
  XOR2_X1 \SubCellInst_LFInst_9_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_9_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_9_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_9_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_1_U12  ( .A1(StateRegOutput[37]), .A2(
        \SubCellInst_LFInst_9_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_1_U11  ( .A1(StateRegOutput[39]), .A2(
        \SubCellInst_LFInst_9_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_9_LFInst_1_U10  ( .A1(StateRegOutput[36]), .A2(
        StateRegOutput[38]), .ZN(\SubCellInst_LFInst_9_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_1_U9  ( .A1(StateRegOutput[39]), .A2(
        \SubCellInst_LFInst_9_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_1_U8  ( .A1(
        \SubCellInst_LFInst_9_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_9_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_1_U7  ( .A1(StateRegOutput[36]), .A2(
        StateRegOutput[38]), .ZN(\SubCellInst_LFInst_9_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_9_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_9_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_1_U5  ( .A1(StateRegOutput[36]), .A2(
        StateRegOutput[37]), .ZN(\SubCellInst_LFInst_9_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_9_LFInst_1_U4  ( .A(StateRegOutput[38]), .ZN(
        \SubCellInst_LFInst_9_LFInst_1_n11 ) );
  NAND2_X2 \SubCellInst_LFInst_9_LFInst_1_U3  ( .A1(
        \SubCellInst_LFInst_9_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_9_LFInst_1_n17 ), .ZN(\Red_MCInst_MC1_v1_2 [1]) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_9_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_9_LFInst_2_n21 ), .ZN(\MCInst_MC1_v1_3 [3]) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U10  ( .A1(StateRegOutput[38]), .A2(
        \SubCellInst_LFInst_9_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_2_U9  ( .A1(StateRegOutput[37]), .A2(
        \SubCellInst_LFInst_9_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_9_LFInst_2_U8  ( .A(StateRegOutput[39]), .ZN(
        \SubCellInst_LFInst_9_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_9_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_9_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_9_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_9_LFInst_2_n16 ), .B(StateRegOutput[38]), .Z(
        \SubCellInst_LFInst_9_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U5  ( .A1(StateRegOutput[36]), .A2(
        StateRegOutput[37]), .ZN(\SubCellInst_LFInst_9_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_9_LFInst_2_n15 ), .A2(StateRegOutput[39]), .ZN(
        \SubCellInst_LFInst_9_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_9_LFInst_2_U3  ( .A(StateRegOutput[36]), .B(
        StateRegOutput[37]), .ZN(\SubCellInst_LFInst_9_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_9_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_9_LFInst_3_n15 ), .ZN(\Red_MCInst_MC1_v1_1 [2]) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_3_U8  ( .A1(StateRegOutput[37]), .A2(
        \SubCellInst_LFInst_9_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_9_LFInst_3_U7  ( .A(StateRegOutput[39]), .B(
        StateRegOutput[38]), .Z(\SubCellInst_LFInst_9_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_9_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_9_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_3_U5  ( .A1(StateRegOutput[36]), .A2(
        StateRegOutput[38]), .ZN(\SubCellInst_LFInst_9_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_9_LFInst_3_U4  ( .A(StateRegOutput[36]), .B(
        \SubCellInst_LFInst_9_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_9_LFInst_3_U3  ( .A1(StateRegOutput[39]), .A2(
        StateRegOutput[37]), .ZN(\SubCellInst_LFInst_9_LFInst_3_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_0_U7  ( .A1(AddConstOutput[18]), .A2(
        \SubCellInst_LFInst_10_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_10_LFInst_0_U6  ( .A(AddConstOutput[17]), .ZN(
        \SubCellInst_LFInst_10_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_10_LFInst_0_U5  ( .A(AddConstOutput[16]), .B(
        AddConstOutput[19]), .Z(\SubCellInst_LFInst_10_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_10_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_10_LFInst_0_n10 ), .ZN(\MCInst_MC0_v1_0 [0]) );
  XOR2_X1 \SubCellInst_LFInst_10_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_10_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_10_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_10_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_1_U12  ( .A1(AddConstOutput[17]), 
        .A2(\SubCellInst_LFInst_10_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_1_U11  ( .A1(AddConstOutput[19]), .A2(
        \SubCellInst_LFInst_10_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_10_LFInst_1_U10  ( .A1(AddConstOutput[16]), .A2(
        AddConstOutput[18]), .ZN(\SubCellInst_LFInst_10_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_1_U9  ( .A1(AddConstOutput[19]), .A2(
        \SubCellInst_LFInst_10_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_1_U8  ( .A1(
        \SubCellInst_LFInst_10_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_10_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_1_U7  ( .A1(AddConstOutput[16]), .A2(
        AddConstOutput[18]), .ZN(\SubCellInst_LFInst_10_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_10_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_10_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_1_U5  ( .A1(AddConstOutput[16]), .A2(
        AddConstOutput[17]), .ZN(\SubCellInst_LFInst_10_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_10_LFInst_1_U4  ( .A(AddConstOutput[18]), .ZN(
        \SubCellInst_LFInst_10_LFInst_1_n11 ) );
  NAND2_X2 \SubCellInst_LFInst_10_LFInst_1_U3  ( .A1(
        \SubCellInst_LFInst_10_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_10_LFInst_1_n17 ), .ZN(\Red_MCInst_MC0_v1_2 [1])
         );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_10_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_10_LFInst_2_n21 ), .ZN(\MCInst_MC0_v1_3 [3]) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U10  ( .A1(AddConstOutput[18]), 
        .A2(\SubCellInst_LFInst_10_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_2_U9  ( .A1(AddConstOutput[17]), .A2(
        \SubCellInst_LFInst_10_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_10_LFInst_2_U8  ( .A(AddConstOutput[19]), .ZN(
        \SubCellInst_LFInst_10_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_10_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_10_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_10_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_10_LFInst_2_n16 ), .B(AddConstOutput[18]), .Z(
        \SubCellInst_LFInst_10_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U5  ( .A1(AddConstOutput[16]), .A2(
        AddConstOutput[17]), .ZN(\SubCellInst_LFInst_10_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_10_LFInst_2_n15 ), .A2(AddConstOutput[19]), .ZN(
        \SubCellInst_LFInst_10_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_10_LFInst_2_U3  ( .A(AddConstOutput[16]), .B(
        AddConstOutput[17]), .ZN(\SubCellInst_LFInst_10_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_10_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_10_LFInst_3_n15 ), .ZN(\Red_MCInst_MC0_v1_1 [2])
         );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_3_U8  ( .A1(AddConstOutput[17]), .A2(
        \SubCellInst_LFInst_10_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_10_LFInst_3_U7  ( .A(AddConstOutput[19]), .B(
        AddConstOutput[18]), .Z(\SubCellInst_LFInst_10_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_10_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_10_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_3_U5  ( .A1(AddConstOutput[16]), .A2(
        AddConstOutput[18]), .ZN(\SubCellInst_LFInst_10_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_10_LFInst_3_U4  ( .A(AddConstOutput[16]), .B(
        \SubCellInst_LFInst_10_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_10_LFInst_3_U3  ( .A1(AddConstOutput[19]), .A2(
        AddConstOutput[17]), .ZN(\SubCellInst_LFInst_10_LFInst_3_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_0_U7  ( .A1(AddConstOutput[22]), .A2(
        \SubCellInst_LFInst_11_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_11_LFInst_0_U6  ( .A(AddConstOutput[21]), .ZN(
        \SubCellInst_LFInst_11_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_11_LFInst_0_U5  ( .A(AddConstOutput[20]), .B(
        AddConstOutput[23]), .Z(\SubCellInst_LFInst_11_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_11_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_11_LFInst_0_n10 ), .ZN(\MCInst_MC3_v1_0 [0]) );
  XOR2_X1 \SubCellInst_LFInst_11_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_11_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_11_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_11_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_1_U12  ( .A1(AddConstOutput[21]), 
        .A2(\SubCellInst_LFInst_11_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_1_U11  ( .A1(AddConstOutput[23]), .A2(
        \SubCellInst_LFInst_11_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_11_LFInst_1_U10  ( .A1(AddConstOutput[20]), .A2(
        AddConstOutput[22]), .ZN(\SubCellInst_LFInst_11_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_1_U9  ( .A1(AddConstOutput[23]), .A2(
        \SubCellInst_LFInst_11_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_1_U8  ( .A1(
        \SubCellInst_LFInst_11_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_11_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_1_U7  ( .A1(AddConstOutput[20]), .A2(
        AddConstOutput[22]), .ZN(\SubCellInst_LFInst_11_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_11_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_11_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_1_U5  ( .A1(AddConstOutput[20]), .A2(
        AddConstOutput[21]), .ZN(\SubCellInst_LFInst_11_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_11_LFInst_1_U4  ( .A(AddConstOutput[22]), .ZN(
        \SubCellInst_LFInst_11_LFInst_1_n11 ) );
  NAND2_X2 \SubCellInst_LFInst_11_LFInst_1_U3  ( .A1(
        \SubCellInst_LFInst_11_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_11_LFInst_1_n17 ), .ZN(\Red_MCInst_MC3_v1_2 [1])
         );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_11_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_11_LFInst_2_n21 ), .ZN(\MCInst_MC3_v1_3 [3]) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U10  ( .A1(AddConstOutput[22]), 
        .A2(\SubCellInst_LFInst_11_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_2_U9  ( .A1(AddConstOutput[21]), .A2(
        \SubCellInst_LFInst_11_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_11_LFInst_2_U8  ( .A(AddConstOutput[23]), .ZN(
        \SubCellInst_LFInst_11_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_11_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_11_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_11_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_11_LFInst_2_n16 ), .B(AddConstOutput[22]), .Z(
        \SubCellInst_LFInst_11_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U5  ( .A1(AddConstOutput[20]), .A2(
        AddConstOutput[21]), .ZN(\SubCellInst_LFInst_11_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_11_LFInst_2_n15 ), .A2(AddConstOutput[23]), .ZN(
        \SubCellInst_LFInst_11_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_11_LFInst_2_U3  ( .A(AddConstOutput[20]), .B(
        AddConstOutput[21]), .ZN(\SubCellInst_LFInst_11_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_11_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_11_LFInst_3_n15 ), .ZN(\Red_MCInst_MC3_v1_1 [2])
         );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_3_U8  ( .A1(AddConstOutput[21]), .A2(
        \SubCellInst_LFInst_11_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_11_LFInst_3_U7  ( .A(AddConstOutput[23]), .B(
        AddConstOutput[22]), .Z(\SubCellInst_LFInst_11_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_11_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_11_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_3_U5  ( .A1(AddConstOutput[20]), .A2(
        AddConstOutput[22]), .ZN(\SubCellInst_LFInst_11_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_11_LFInst_3_U4  ( .A(AddConstOutput[20]), .B(
        \SubCellInst_LFInst_11_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_11_LFInst_3_U3  ( .A1(AddConstOutput[23]), .A2(
        AddConstOutput[21]), .ZN(\SubCellInst_LFInst_11_LFInst_3_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_0_U7  ( .A1(StateRegOutput[50]), .A2(
        \SubCellInst_LFInst_12_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_12_LFInst_0_U6  ( .A(StateRegOutput[49]), .ZN(
        \SubCellInst_LFInst_12_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_12_LFInst_0_U5  ( .A(StateRegOutput[48]), .B(
        StateRegOutput[51]), .Z(\SubCellInst_LFInst_12_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_12_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_12_LFInst_0_n10 ), .ZN(\Red_MCInst_MC3_v0_0 [0])
         );
  XOR2_X1 \SubCellInst_LFInst_12_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_12_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_12_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_12_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_12_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_12_LFInst_1_n17 ), .ZN(\Red_MCInst_MC3_v0_2 [2])
         );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U11  ( .A1(StateRegOutput[49]), 
        .A2(\SubCellInst_LFInst_12_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_1_U10  ( .A1(StateRegOutput[51]), .A2(
        \SubCellInst_LFInst_12_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_12_LFInst_1_U9  ( .A1(StateRegOutput[48]), .A2(
        StateRegOutput[50]), .ZN(\SubCellInst_LFInst_12_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U8  ( .A1(StateRegOutput[51]), .A2(
        \SubCellInst_LFInst_12_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_12_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_12_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U6  ( .A1(StateRegOutput[48]), .A2(
        StateRegOutput[50]), .ZN(\SubCellInst_LFInst_12_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_12_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_12_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U4  ( .A1(StateRegOutput[48]), .A2(
        StateRegOutput[49]), .ZN(\SubCellInst_LFInst_12_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_12_LFInst_1_U3  ( .A(StateRegOutput[50]), .ZN(
        \SubCellInst_LFInst_12_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_12_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_12_LFInst_2_n21 ), .ZN(\MCInst_MC3_v0_3 [3]) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U10  ( .A1(StateRegOutput[50]), 
        .A2(\SubCellInst_LFInst_12_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_2_U9  ( .A1(StateRegOutput[49]), .A2(
        \SubCellInst_LFInst_12_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_12_LFInst_2_U8  ( .A(StateRegOutput[51]), .ZN(
        \SubCellInst_LFInst_12_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_12_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_12_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_12_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_12_LFInst_2_n16 ), .B(StateRegOutput[50]), .Z(
        \SubCellInst_LFInst_12_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U5  ( .A1(StateRegOutput[48]), .A2(
        StateRegOutput[49]), .ZN(\SubCellInst_LFInst_12_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_12_LFInst_2_n15 ), .A2(StateRegOutput[51]), .ZN(
        \SubCellInst_LFInst_12_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_12_LFInst_2_U3  ( .A(StateRegOutput[48]), .B(
        StateRegOutput[49]), .ZN(\SubCellInst_LFInst_12_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_12_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_12_LFInst_3_n15 ), .ZN(\Red_MCInst_MC3_v0_1 [0])
         );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_3_U8  ( .A1(StateRegOutput[49]), .A2(
        \SubCellInst_LFInst_12_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_12_LFInst_3_U7  ( .A(StateRegOutput[51]), .B(
        StateRegOutput[50]), .Z(\SubCellInst_LFInst_12_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_12_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_12_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_3_U5  ( .A1(StateRegOutput[48]), .A2(
        StateRegOutput[50]), .ZN(\SubCellInst_LFInst_12_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_12_LFInst_3_U4  ( .A(StateRegOutput[48]), .B(
        \SubCellInst_LFInst_12_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_12_LFInst_3_U3  ( .A1(StateRegOutput[51]), .A2(
        StateRegOutput[49]), .ZN(\SubCellInst_LFInst_12_LFInst_3_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_0_U7  ( .A1(StateRegOutput[54]), .A2(
        \SubCellInst_LFInst_13_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_13_LFInst_0_U6  ( .A(StateRegOutput[53]), .ZN(
        \SubCellInst_LFInst_13_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_13_LFInst_0_U5  ( .A(StateRegOutput[52]), .B(
        StateRegOutput[55]), .Z(\SubCellInst_LFInst_13_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_13_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_13_LFInst_0_n10 ), .ZN(\Red_MCInst_MC2_v0_0 [0])
         );
  XOR2_X1 \SubCellInst_LFInst_13_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_13_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_13_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_13_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_13_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_13_LFInst_1_n17 ), .ZN(\Red_MCInst_MC2_v0_2 [2])
         );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U11  ( .A1(StateRegOutput[53]), 
        .A2(\SubCellInst_LFInst_13_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_1_U10  ( .A1(StateRegOutput[55]), .A2(
        \SubCellInst_LFInst_13_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_13_LFInst_1_U9  ( .A1(StateRegOutput[52]), .A2(
        StateRegOutput[54]), .ZN(\SubCellInst_LFInst_13_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U8  ( .A1(StateRegOutput[55]), .A2(
        \SubCellInst_LFInst_13_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_13_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_13_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U6  ( .A1(StateRegOutput[52]), .A2(
        StateRegOutput[54]), .ZN(\SubCellInst_LFInst_13_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_13_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_13_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U4  ( .A1(StateRegOutput[52]), .A2(
        StateRegOutput[53]), .ZN(\SubCellInst_LFInst_13_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_13_LFInst_1_U3  ( .A(StateRegOutput[54]), .ZN(
        \SubCellInst_LFInst_13_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_13_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_13_LFInst_2_n21 ), .ZN(\MCInst_MC2_v0_3 [3]) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U10  ( .A1(StateRegOutput[54]), 
        .A2(\SubCellInst_LFInst_13_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_2_U9  ( .A1(StateRegOutput[53]), .A2(
        \SubCellInst_LFInst_13_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_13_LFInst_2_U8  ( .A(StateRegOutput[55]), .ZN(
        \SubCellInst_LFInst_13_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_13_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_13_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_13_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_13_LFInst_2_n16 ), .B(StateRegOutput[54]), .Z(
        \SubCellInst_LFInst_13_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U5  ( .A1(StateRegOutput[52]), .A2(
        StateRegOutput[53]), .ZN(\SubCellInst_LFInst_13_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_13_LFInst_2_n15 ), .A2(StateRegOutput[55]), .ZN(
        \SubCellInst_LFInst_13_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_13_LFInst_2_U3  ( .A(StateRegOutput[52]), .B(
        StateRegOutput[53]), .ZN(\SubCellInst_LFInst_13_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_13_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_13_LFInst_3_n15 ), .ZN(\Red_MCInst_MC2_v0_1 [0])
         );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_3_U8  ( .A1(StateRegOutput[53]), .A2(
        \SubCellInst_LFInst_13_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_13_LFInst_3_U7  ( .A(StateRegOutput[55]), .B(
        StateRegOutput[54]), .Z(\SubCellInst_LFInst_13_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_13_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_13_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_3_U5  ( .A1(StateRegOutput[52]), .A2(
        StateRegOutput[54]), .ZN(\SubCellInst_LFInst_13_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_13_LFInst_3_U4  ( .A(StateRegOutput[52]), .B(
        \SubCellInst_LFInst_13_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_13_LFInst_3_U3  ( .A1(StateRegOutput[55]), .A2(
        StateRegOutput[53]), .ZN(\SubCellInst_LFInst_13_LFInst_3_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_0_U7  ( .A1(AddConstOutput[26]), .A2(
        \SubCellInst_LFInst_14_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_14_LFInst_0_U6  ( .A(AddConstOutput[25]), .ZN(
        \SubCellInst_LFInst_14_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_14_LFInst_0_U5  ( .A(AddConstOutput[24]), .B(
        AddConstOutput[27]), .Z(\SubCellInst_LFInst_14_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_14_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_14_LFInst_0_n10 ), .ZN(\Red_MCInst_MC1_v0_0 [0])
         );
  XOR2_X1 \SubCellInst_LFInst_14_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_14_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_14_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_14_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_14_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_14_LFInst_1_n17 ), .ZN(\Red_MCInst_MC1_v0_2 [2])
         );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U11  ( .A1(AddConstOutput[25]), 
        .A2(\SubCellInst_LFInst_14_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_1_U10  ( .A1(AddConstOutput[27]), .A2(
        \SubCellInst_LFInst_14_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_14_LFInst_1_U9  ( .A1(AddConstOutput[24]), .A2(
        AddConstOutput[26]), .ZN(\SubCellInst_LFInst_14_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U8  ( .A1(AddConstOutput[27]), .A2(
        \SubCellInst_LFInst_14_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_14_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_14_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U6  ( .A1(AddConstOutput[24]), .A2(
        AddConstOutput[26]), .ZN(\SubCellInst_LFInst_14_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_14_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_14_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U4  ( .A1(AddConstOutput[24]), .A2(
        AddConstOutput[25]), .ZN(\SubCellInst_LFInst_14_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_14_LFInst_1_U3  ( .A(AddConstOutput[26]), .ZN(
        \SubCellInst_LFInst_14_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_14_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_14_LFInst_2_n21 ), .ZN(\MCInst_MC1_v0_3 [3]) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U10  ( .A1(AddConstOutput[26]), 
        .A2(\SubCellInst_LFInst_14_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_2_U9  ( .A1(AddConstOutput[25]), .A2(
        \SubCellInst_LFInst_14_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_14_LFInst_2_U8  ( .A(AddConstOutput[27]), .ZN(
        \SubCellInst_LFInst_14_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_14_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_14_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_14_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_14_LFInst_2_n16 ), .B(AddConstOutput[26]), .Z(
        \SubCellInst_LFInst_14_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U5  ( .A1(AddConstOutput[24]), .A2(
        AddConstOutput[25]), .ZN(\SubCellInst_LFInst_14_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_14_LFInst_2_n15 ), .A2(AddConstOutput[27]), .ZN(
        \SubCellInst_LFInst_14_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_14_LFInst_2_U3  ( .A(AddConstOutput[24]), .B(
        AddConstOutput[25]), .ZN(\SubCellInst_LFInst_14_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_14_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_14_LFInst_3_n15 ), .ZN(\Red_MCInst_MC1_v0_1 [0])
         );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_3_U8  ( .A1(AddConstOutput[25]), .A2(
        \SubCellInst_LFInst_14_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_14_LFInst_3_U7  ( .A(AddConstOutput[27]), .B(
        AddConstOutput[26]), .Z(\SubCellInst_LFInst_14_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_14_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_14_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_3_U5  ( .A1(AddConstOutput[24]), .A2(
        AddConstOutput[26]), .ZN(\SubCellInst_LFInst_14_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_14_LFInst_3_U4  ( .A(AddConstOutput[24]), .B(
        \SubCellInst_LFInst_14_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_14_LFInst_3_U3  ( .A1(AddConstOutput[27]), .A2(
        AddConstOutput[25]), .ZN(\SubCellInst_LFInst_14_LFInst_3_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_0_U7  ( .A1(AddConstOutput[30]), .A2(
        \SubCellInst_LFInst_15_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_15_LFInst_0_U6  ( .A(AddConstOutput[29]), .ZN(
        \SubCellInst_LFInst_15_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_15_LFInst_0_U5  ( .A(AddConstOutput[28]), .B(
        AddConstOutput[31]), .Z(\SubCellInst_LFInst_15_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_15_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_15_LFInst_0_n10 ), .ZN(\Red_MCInst_MC0_v0_0 [0])
         );
  XOR2_X1 \SubCellInst_LFInst_15_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_15_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_15_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_15_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_15_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_15_LFInst_1_n17 ), .ZN(\Red_MCInst_MC0_v0_2 [2])
         );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U11  ( .A1(AddConstOutput[29]), 
        .A2(\SubCellInst_LFInst_15_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_1_U10  ( .A1(AddConstOutput[31]), .A2(
        \SubCellInst_LFInst_15_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_15_LFInst_1_U9  ( .A1(AddConstOutput[28]), .A2(
        AddConstOutput[30]), .ZN(\SubCellInst_LFInst_15_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U8  ( .A1(AddConstOutput[31]), .A2(
        \SubCellInst_LFInst_15_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_15_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_15_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U6  ( .A1(AddConstOutput[28]), .A2(
        AddConstOutput[30]), .ZN(\SubCellInst_LFInst_15_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_15_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_15_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U4  ( .A1(AddConstOutput[28]), .A2(
        AddConstOutput[29]), .ZN(\SubCellInst_LFInst_15_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_15_LFInst_1_U3  ( .A(AddConstOutput[30]), .ZN(
        \SubCellInst_LFInst_15_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_15_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_15_LFInst_2_n21 ), .ZN(\MCInst_MC0_v0_3 [3]) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U10  ( .A1(AddConstOutput[30]), 
        .A2(\SubCellInst_LFInst_15_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_2_U9  ( .A1(AddConstOutput[29]), .A2(
        \SubCellInst_LFInst_15_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_15_LFInst_2_U8  ( .A(AddConstOutput[31]), .ZN(
        \SubCellInst_LFInst_15_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_15_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_15_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_15_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_15_LFInst_2_n16 ), .B(AddConstOutput[30]), .Z(
        \SubCellInst_LFInst_15_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U5  ( .A1(AddConstOutput[28]), .A2(
        AddConstOutput[29]), .ZN(\SubCellInst_LFInst_15_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_15_LFInst_2_n15 ), .A2(AddConstOutput[31]), .ZN(
        \SubCellInst_LFInst_15_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_15_LFInst_2_U3  ( .A(AddConstOutput[28]), .B(
        AddConstOutput[29]), .ZN(\SubCellInst_LFInst_15_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_15_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_15_LFInst_3_n15 ), .ZN(\Red_MCInst_MC0_v0_1 [0])
         );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_3_U8  ( .A1(AddConstOutput[29]), .A2(
        \SubCellInst_LFInst_15_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_15_LFInst_3_U7  ( .A(AddConstOutput[31]), .B(
        AddConstOutput[30]), .Z(\SubCellInst_LFInst_15_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_15_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_15_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_3_U5  ( .A1(AddConstOutput[28]), .A2(
        AddConstOutput[30]), .ZN(\SubCellInst_LFInst_15_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_15_LFInst_3_U4  ( .A(AddConstOutput[28]), .B(
        \SubCellInst_LFInst_15_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_15_LFInst_3_U3  ( .A1(AddConstOutput[31]), .A2(
        AddConstOutput[29]), .ZN(\SubCellInst_LFInst_15_LFInst_3_n11 ) );
  XNOR2_X1 \MCInst_MC0_v0_2Inst_0_U4  ( .A(\MCInst_MC0_v0_2Inst_0_n2 ), .B(
        \Red_MCInst_MC0_v0_2 [2]), .ZN(\MCInst_MC0_v0_2 [0]) );
  XNOR2_X1 \MCInst_MC0_v0_2Inst_0_U3  ( .A(\Red_MCInst_MC0_v0_1 [0]), .B(
        \Red_MCInst_MC0_v0_0 [0]), .ZN(\MCInst_MC0_v0_2Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC0_v1_1Inst_0_U3  ( .A(\MCInst_MC0_v1_3 [3]), .B(
        \Red_MCInst_MC0_v1_1 [2]), .Z(\MCInst_MC0_v1_1 [0]) );
  XNOR2_X1 \MCInst_MC0_v1_2Inst_0_U4  ( .A(\MCInst_MC0_v1_2Inst_0_n2 ), .B(
        \MCInst_MC0_v1_3 [3]), .ZN(\MCInst_MC0_v1_2 [0]) );
  XNOR2_X1 \MCInst_MC0_v1_2Inst_0_U3  ( .A(\Red_MCInst_MC0_v1_1 [2]), .B(
        \Red_MCInst_MC0_v1_2 [1]), .ZN(\MCInst_MC0_v1_2Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC0_v2_1Inst_0_U3  ( .A(\Red_MCInst_MC0_v2_1 [1]), .B(
        \MCInst_MC0_v2_0 [3]), .Z(\MCInst_MC0_v2_1 [0]) );
  XOR2_X1 \MCInst_MC0_v2_2Inst_0_U3  ( .A(\MCInst_MC0_v2_0 [2]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\MCInst_MC0_v2_2 [0]) );
  XNOR2_X1 \MCInst_MC0_v2_3Inst_0_U5  ( .A(\MCInst_MC0_v2_3Inst_0_n4 ), .B(
        \MCInst_MC0_v2_3Inst_0_n3 ), .ZN(\MCInst_MC0_v2_3 [0]) );
  XNOR2_X1 \MCInst_MC0_v2_3Inst_0_U4  ( .A(\MCInst_MC0_v2_0 [2]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\MCInst_MC0_v2_3Inst_0_n3 ) );
  XOR2_X1 \MCInst_MC0_v2_3Inst_0_U3  ( .A(\MCInst_MC0_v2_0 [3]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\MCInst_MC0_v2_3Inst_0_n4 ) );
  XOR2_X1 \MCInst_MC0_v3_1Inst_0_U3  ( .A(\MCInst_MC0_v3_0 [3]), .B(
        \Red_MCInst_MC0_v3_1 [2]), .Z(\MCInst_MC0_v3_1 [0]) );
  XOR2_X1 \MCInst_MC0_v3_2Inst_0_U3  ( .A(\MCInst_MC0_v3_2 [3]), .B(
        \Red_MCInst_MC0_v3_3 [2]), .Z(\MCInst_MC0_v3_2 [0]) );
  XNOR2_X1 \MCInst_MC0_v3_3Inst_0_U4  ( .A(\MCInst_MC0_v3_3Inst_0_n2 ), .B(
        \Red_MCInst_MC0_v3_3 [2]), .ZN(\MCInst_MC0_v3_3 [0]) );
  XNOR2_X1 \MCInst_MC0_v3_3Inst_0_U3  ( .A(\Red_MCInst_MC0_v3_1 [2]), .B(
        \MCInst_MC0_v3_2 [3]), .ZN(\MCInst_MC0_v3_3Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC0_v0_0Inst_1_U3  ( .A(\MCInst_MC0_v0_3 [3]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\MCInst_MC0_v0_0 [1]) );
  XOR2_X1 \MCInst_MC0_v0_1Inst_1_U3  ( .A(\Red_MCInst_MC0_v0_2 [2]), .B(
        \MCInst_MC0_v0_3 [3]), .Z(\MCInst_MC0_v0_1 [1]) );
  XNOR2_X1 \MCInst_MC0_v0_2Inst_1_U4  ( .A(\MCInst_MC0_v0_2Inst_1_n2 ), .B(
        \MCInst_MC0_v0_3 [3]), .ZN(\MCInst_MC0_v0_2 [1]) );
  XNOR2_X1 \MCInst_MC0_v0_2Inst_1_U3  ( .A(\Red_MCInst_MC0_v0_1 [0]), .B(
        \Red_MCInst_MC0_v0_0 [0]), .ZN(\MCInst_MC0_v0_2Inst_1_n2 ) );
  XOR2_X1 \MCInst_MC0_v0_3Inst_1_U3  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\MCInst_MC0_v0_3 [1]) );
  XOR2_X1 \MCInst_MC0_v1_1Inst_1_U3  ( .A(\MCInst_MC0_v1_0 [0]), .B(
        \MCInst_MC0_v1_3 [3]), .Z(\MCInst_MC0_v1_1 [1]) );
  XOR2_X1 \MCInst_MC0_v1_2Inst_1_U3  ( .A(\MCInst_MC0_v1_0 [0]), .B(
        \Red_MCInst_MC0_v1_2 [1]), .Z(\MCInst_MC0_v1_2 [1]) );
  XOR2_X1 \MCInst_MC0_v1_3Inst_1_U3  ( .A(\MCInst_MC0_v1_0 [0]), .B(
        \Red_MCInst_MC0_v1_1 [2]), .Z(\MCInst_MC0_v1_3 [1]) );
  XOR2_X1 \MCInst_MC0_v2_0Inst_1_U3  ( .A(\Red_MCInst_MC0_v2_1 [1]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\MCInst_MC0_v2_0 [1]) );
  XNOR2_X1 \MCInst_MC0_v2_1Inst_1_U4  ( .A(\MCInst_MC0_v2_1Inst_1_n2 ), .B(
        \MCInst_MC0_v2_0 [3]), .ZN(\MCInst_MC0_v2_1 [1]) );
  XNOR2_X1 \MCInst_MC0_v2_1Inst_1_U3  ( .A(\Red_MCInst_MC0_v2_2 [1]), .B(
        \MCInst_MC0_v2_0 [2]), .ZN(\MCInst_MC0_v2_1Inst_1_n2 ) );
  XNOR2_X1 \MCInst_MC0_v2_2Inst_1_U5  ( .A(\MCInst_MC0_v2_2Inst_1_n4 ), .B(
        \MCInst_MC0_v2_2Inst_1_n3 ), .ZN(\MCInst_MC0_v2_2 [1]) );
  XNOR2_X1 \MCInst_MC0_v2_2Inst_1_U4  ( .A(\MCInst_MC0_v2_0 [2]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\MCInst_MC0_v2_2Inst_1_n3 ) );
  XOR2_X1 \MCInst_MC0_v2_2Inst_1_U3  ( .A(\MCInst_MC0_v2_0 [3]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\MCInst_MC0_v2_2Inst_1_n4 ) );
  XOR2_X1 \MCInst_MC0_v3_0Inst_1_U3  ( .A(\MCInst_MC0_v3_2 [3]), .B(
        \Red_MCInst_MC0_v3_1 [2]), .Z(\MCInst_MC0_v3_0 [1]) );
  XOR2_X1 \MCInst_MC0_v3_1Inst_1_U3  ( .A(\MCInst_MC0_v3_2 [3]), .B(
        \MCInst_MC0_v3_0 [3]), .Z(\MCInst_MC0_v3_1 [1]) );
  XNOR2_X1 \MCInst_MC0_v3_3Inst_1_U4  ( .A(\MCInst_MC0_v3_3Inst_1_n2 ), .B(
        \MCInst_MC0_v3_0 [3]), .ZN(\MCInst_MC0_v3_3 [1]) );
  XNOR2_X1 \MCInst_MC0_v3_3Inst_1_U3  ( .A(\Red_MCInst_MC0_v3_1 [2]), .B(
        \MCInst_MC0_v3_2 [3]), .ZN(\MCInst_MC0_v3_3Inst_1_n2 ) );
  XOR2_X1 \MCInst_MC0_v0_0Inst_2_U3  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\MCInst_MC0_v0_0 [2]) );
  XOR2_X1 \MCInst_MC0_v0_1Inst_2_U3  ( .A(\MCInst_MC0_v0_3 [3]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\MCInst_MC0_v0_1 [2]) );
  XOR2_X1 \MCInst_MC0_v0_2Inst_2_U3  ( .A(\Red_MCInst_MC0_v0_2 [2]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\MCInst_MC0_v0_2 [2]) );
  XNOR2_X1 \MCInst_MC0_v1_1Inst_2_U4  ( .A(\MCInst_MC0_v1_1Inst_2_n2 ), .B(
        \Red_MCInst_MC0_v1_2 [1]), .ZN(\MCInst_MC0_v1_1 [2]) );
  XNOR2_X1 \MCInst_MC0_v1_1Inst_2_U3  ( .A(\Red_MCInst_MC0_v1_1 [2]), .B(
        \MCInst_MC0_v1_0 [0]), .ZN(\MCInst_MC0_v1_1Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC0_v1_2Inst_2_U4  ( .A(\MCInst_MC0_v1_2Inst_2_n2 ), .B(
        \Red_MCInst_MC0_v1_2 [1]), .ZN(\MCInst_MC0_v1_2 [2]) );
  XNOR2_X1 \MCInst_MC0_v1_2Inst_2_U3  ( .A(\MCInst_MC0_v1_3 [3]), .B(
        \MCInst_MC0_v1_0 [0]), .ZN(\MCInst_MC0_v1_2Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC0_v2_1Inst_2_U4  ( .A(\MCInst_MC0_v2_1Inst_2_n2 ), .B(
        \MCInst_MC0_v2_0 [3]), .ZN(\MCInst_MC0_v2_1 [2]) );
  XNOR2_X1 \MCInst_MC0_v2_1Inst_2_U3  ( .A(\Red_MCInst_MC0_v2_2 [1]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\MCInst_MC0_v2_1Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC0_v2_2Inst_2_U4  ( .A(\MCInst_MC0_v2_2Inst_2_n2 ), .B(
        \MCInst_MC0_v2_0 [3]), .ZN(\MCInst_MC0_v2_2 [2]) );
  XNOR2_X1 \MCInst_MC0_v2_2Inst_2_U3  ( .A(\Red_MCInst_MC0_v2_2 [1]), .B(
        \MCInst_MC0_v2_0 [2]), .ZN(\MCInst_MC0_v2_2Inst_2_n2 ) );
  XOR2_X1 \MCInst_MC0_v2_3Inst_2_U3  ( .A(\Red_MCInst_MC0_v2_1 [1]), .B(
        \MCInst_MC0_v2_0 [2]), .Z(\MCInst_MC0_v2_3 [2]) );
  XNOR2_X1 \MCInst_MC0_v3_1Inst_2_U4  ( .A(\MCInst_MC0_v3_1Inst_2_n2 ), .B(
        \Red_MCInst_MC0_v3_3 [2]), .ZN(\MCInst_MC0_v3_1 [2]) );
  XNOR2_X1 \MCInst_MC0_v3_1Inst_2_U3  ( .A(\Red_MCInst_MC0_v3_1 [2]), .B(
        \MCInst_MC0_v3_2 [3]), .ZN(\MCInst_MC0_v3_1Inst_2_n2 ) );
  XOR2_X1 \MCInst_MC0_v3_3Inst_2_U3  ( .A(\Red_MCInst_MC0_v3_3 [2]), .B(
        \Red_MCInst_MC0_v3_1 [2]), .Z(\MCInst_MC0_v3_3 [2]) );
  XOR2_X1 \MCInst_MC0_v0_1Inst_3_U3  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\MCInst_MC0_v0_1 [3]) );
  XOR2_X1 \MCInst_MC0_v0_2Inst_3_U3  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(
        \MCInst_MC0_v0_3 [3]), .Z(\MCInst_MC0_v0_2 [3]) );
  XOR2_X1 \MCInst_MC0_v1_1Inst_3_U3  ( .A(\Red_MCInst_MC0_v1_2 [1]), .B(
        \MCInst_MC0_v1_3 [3]), .Z(\MCInst_MC0_v1_1 [3]) );
  XNOR2_X1 \MCInst_MC0_v1_2Inst_3_U5  ( .A(\MCInst_MC0_v1_2Inst_3_n4 ), .B(
        \MCInst_MC0_v1_2Inst_3_n3 ), .ZN(\MCInst_MC0_v1_2 [3]) );
  XNOR2_X1 \MCInst_MC0_v1_2Inst_3_U4  ( .A(\Red_MCInst_MC0_v1_2 [1]), .B(
        \MCInst_MC0_v1_0 [0]), .ZN(\MCInst_MC0_v1_2Inst_3_n3 ) );
  XOR2_X1 \MCInst_MC0_v1_2Inst_3_U3  ( .A(\MCInst_MC0_v1_3 [3]), .B(
        \Red_MCInst_MC0_v1_1 [2]), .Z(\MCInst_MC0_v1_2Inst_3_n4 ) );
  XOR2_X1 \MCInst_MC0_v2_1Inst_3_U3  ( .A(\MCInst_MC0_v2_0 [2]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\MCInst_MC0_v2_1 [3]) );
  XNOR2_X1 \MCInst_MC0_v2_2Inst_3_U4  ( .A(\MCInst_MC0_v2_2Inst_3_n2 ), .B(
        \MCInst_MC0_v2_0 [3]), .ZN(\MCInst_MC0_v2_2 [3]) );
  XNOR2_X1 \MCInst_MC0_v2_2Inst_3_U3  ( .A(\Red_MCInst_MC0_v2_2 [1]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\MCInst_MC0_v2_2Inst_3_n2 ) );
  XNOR2_X1 \MCInst_MC0_v2_3Inst_3_U4  ( .A(\MCInst_MC0_v2_3Inst_3_n2 ), .B(
        \MCInst_MC0_v2_0 [2]), .ZN(\MCInst_MC0_v2_3 [3]) );
  XNOR2_X1 \MCInst_MC0_v2_3Inst_3_U3  ( .A(\MCInst_MC0_v2_0 [3]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\MCInst_MC0_v2_3Inst_3_n2 ) );
  XOR2_X1 \MCInst_MC0_v3_1Inst_3_U3  ( .A(\Red_MCInst_MC0_v3_3 [2]), .B(
        \MCInst_MC0_v3_0 [3]), .Z(\MCInst_MC0_v3_1 [3]) );
  XOR2_X1 \MCInst_MC0_v3_3Inst_3_U3  ( .A(\MCInst_MC0_v3_2 [3]), .B(
        \MCInst_MC0_v3_0 [3]), .Z(\MCInst_MC0_v3_3 [3]) );
  XNOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC0_r0Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC0_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[60]) );
  XNOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_0_U2  ( .A(\Red_MCInst_MC0_v3_1 [2]), 
        .B(\Red_MCInst_MC0_v2_2 [1]), .ZN(\MCInst_MC0_r0Inst_XORInst_0_0_n4 )
         );
  XOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_0_U1  ( .A(\MCInst_MC0_v0_3 [3]), .B(
        \MCInst_MC0_v1_0 [0]), .Z(\MCInst_MC0_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC0_r0Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC0_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[61]) );
  XNOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_1_U2  ( .A(\MCInst_MC0_v3_0 [1]), .B(
        \MCInst_MC0_v2_0 [1]), .ZN(\MCInst_MC0_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_1_U1  ( .A(\MCInst_MC0_v0_0 [1]), .B(
        \Red_MCInst_MC0_v1_2 [1]), .Z(\MCInst_MC0_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC0_r0Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC0_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[62]) );
  XNOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_2_U2  ( .A(\Red_MCInst_MC0_v3_3 [2]), 
        .B(\MCInst_MC0_v2_0 [2]), .ZN(\MCInst_MC0_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_2_U1  ( .A(\MCInst_MC0_v0_0 [2]), .B(
        \MCInst_MC0_v1_3 [3]), .Z(\MCInst_MC0_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC0_r0Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC0_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[63]) );
  XNOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_3_U2  ( .A(\MCInst_MC0_v3_0 [3]), .B(
        \MCInst_MC0_v2_0 [3]), .ZN(\MCInst_MC0_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_3_U1  ( .A(\Red_MCInst_MC0_v0_2 [2]), 
        .B(\Red_MCInst_MC0_v1_1 [2]), .Z(\MCInst_MC0_r0Inst_XORInst_0_3_n5 )
         );
  XNOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC0_r1Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC0_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[44]) );
  XNOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_0_U2  ( .A(\MCInst_MC0_v3_1 [0]), .B(
        \MCInst_MC0_v2_1 [0]), .ZN(\MCInst_MC0_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC0_v0_2 [2]), 
        .B(\MCInst_MC0_v1_1 [0]), .Z(\MCInst_MC0_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC0_r1Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC0_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[45]) );
  XNOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_1_U2  ( .A(\MCInst_MC0_v3_1 [1]), .B(
        \MCInst_MC0_v2_1 [1]), .ZN(\MCInst_MC0_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_1_U1  ( .A(\MCInst_MC0_v0_1 [1]), .B(
        \MCInst_MC0_v1_1 [1]), .Z(\MCInst_MC0_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC0_r1Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC0_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[46]) );
  XNOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_2_U2  ( .A(\MCInst_MC0_v3_1 [2]), .B(
        \MCInst_MC0_v2_1 [2]), .ZN(\MCInst_MC0_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_2_U1  ( .A(\MCInst_MC0_v0_1 [2]), .B(
        \MCInst_MC0_v1_1 [2]), .Z(\MCInst_MC0_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC0_r1Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC0_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[47]) );
  XNOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_3_U2  ( .A(\MCInst_MC0_v3_1 [3]), .B(
        \MCInst_MC0_v2_1 [3]), .ZN(\MCInst_MC0_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_3_U1  ( .A(\MCInst_MC0_v0_1 [3]), .B(
        \MCInst_MC0_v1_1 [3]), .Z(\MCInst_MC0_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC0_r2Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC0_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[28]) );
  XNOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_0_U2  ( .A(\MCInst_MC0_v3_2 [0]), .B(
        \MCInst_MC0_v2_2 [0]), .ZN(\MCInst_MC0_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_0_U1  ( .A(\MCInst_MC0_v0_2 [0]), .B(
        \MCInst_MC0_v1_2 [0]), .Z(\MCInst_MC0_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC0_r2Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC0_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[29]) );
  XNOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_1_U2  ( .A(\MCInst_MC0_v3_0 [3]), .B(
        \MCInst_MC0_v2_2 [1]), .ZN(\MCInst_MC0_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_1_U1  ( .A(\MCInst_MC0_v0_2 [1]), .B(
        \MCInst_MC0_v1_2 [1]), .Z(\MCInst_MC0_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC0_r2Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC0_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[30]) );
  XNOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_2_U2  ( .A(\Red_MCInst_MC0_v3_1 [2]), 
        .B(\MCInst_MC0_v2_2 [2]), .ZN(\MCInst_MC0_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_2_U1  ( .A(\MCInst_MC0_v0_2 [2]), .B(
        \MCInst_MC0_v1_2 [2]), .Z(\MCInst_MC0_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC0_r2Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC0_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[31]) );
  XNOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_3_U2  ( .A(\MCInst_MC0_v3_2 [3]), .B(
        \MCInst_MC0_v2_2 [3]), .ZN(\MCInst_MC0_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_3_U1  ( .A(\MCInst_MC0_v0_2 [3]), .B(
        \MCInst_MC0_v1_2 [3]), .Z(\MCInst_MC0_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC0_r3Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC0_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[12]) );
  XNOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_0_U2  ( .A(\MCInst_MC0_v3_3 [0]), .B(
        \MCInst_MC0_v2_3 [0]), .ZN(\MCInst_MC0_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC0_v0_1 [0]), 
        .B(\Red_MCInst_MC0_v1_1 [2]), .Z(\MCInst_MC0_r3Inst_XORInst_0_0_n5 )
         );
  XNOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC0_r3Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC0_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[13]) );
  XNOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_1_U2  ( .A(\MCInst_MC0_v3_3 [1]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\MCInst_MC0_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_1_U1  ( .A(\MCInst_MC0_v0_3 [1]), .B(
        \MCInst_MC0_v1_3 [1]), .Z(\MCInst_MC0_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC0_r3Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC0_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[14]) );
  XNOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_2_U2  ( .A(\MCInst_MC0_v3_3 [2]), .B(
        \MCInst_MC0_v2_3 [2]), .ZN(\MCInst_MC0_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC0_v0_2 [2]), 
        .B(\Red_MCInst_MC0_v1_2 [1]), .Z(\MCInst_MC0_r3Inst_XORInst_0_2_n5 )
         );
  XNOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC0_r3Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC0_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[15]) );
  XNOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_3_U2  ( .A(\MCInst_MC0_v3_3 [3]), .B(
        \MCInst_MC0_v2_3 [3]), .ZN(\MCInst_MC0_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_3_U1  ( .A(\MCInst_MC0_v0_3 [3]), .B(
        \MCInst_MC0_v1_3 [3]), .Z(\MCInst_MC0_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC1_v0_2Inst_0_U4  ( .A(\MCInst_MC1_v0_2Inst_0_n2 ), .B(
        \Red_MCInst_MC1_v0_2 [2]), .ZN(\MCInst_MC1_v0_2 [0]) );
  XNOR2_X1 \MCInst_MC1_v0_2Inst_0_U3  ( .A(\Red_MCInst_MC1_v0_1 [0]), .B(
        \Red_MCInst_MC1_v0_0 [0]), .ZN(\MCInst_MC1_v0_2Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC1_v1_1Inst_0_U3  ( .A(\MCInst_MC1_v1_3 [3]), .B(
        \Red_MCInst_MC1_v1_1 [2]), .Z(\MCInst_MC1_v1_1 [0]) );
  XNOR2_X1 \MCInst_MC1_v1_2Inst_0_U4  ( .A(\MCInst_MC1_v1_2Inst_0_n2 ), .B(
        \MCInst_MC1_v1_3 [3]), .ZN(\MCInst_MC1_v1_2 [0]) );
  XNOR2_X1 \MCInst_MC1_v1_2Inst_0_U3  ( .A(\Red_MCInst_MC1_v1_1 [2]), .B(
        \Red_MCInst_MC1_v1_2 [1]), .ZN(\MCInst_MC1_v1_2Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC1_v2_1Inst_0_U3  ( .A(\Red_MCInst_MC1_v2_1 [1]), .B(
        \MCInst_MC1_v2_0 [3]), .Z(\MCInst_MC1_v2_1 [0]) );
  XOR2_X1 \MCInst_MC1_v2_2Inst_0_U3  ( .A(\MCInst_MC1_v2_0 [2]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\MCInst_MC1_v2_2 [0]) );
  XNOR2_X1 \MCInst_MC1_v2_3Inst_0_U5  ( .A(\MCInst_MC1_v2_3Inst_0_n4 ), .B(
        \MCInst_MC1_v2_3Inst_0_n3 ), .ZN(\MCInst_MC1_v2_3 [0]) );
  XNOR2_X1 \MCInst_MC1_v2_3Inst_0_U4  ( .A(\MCInst_MC1_v2_0 [2]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\MCInst_MC1_v2_3Inst_0_n3 ) );
  XOR2_X1 \MCInst_MC1_v2_3Inst_0_U3  ( .A(\MCInst_MC1_v2_0 [3]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\MCInst_MC1_v2_3Inst_0_n4 ) );
  XOR2_X1 \MCInst_MC1_v3_1Inst_0_U3  ( .A(\MCInst_MC1_v3_0 [3]), .B(
        \Red_MCInst_MC1_v3_1 [2]), .Z(\MCInst_MC1_v3_1 [0]) );
  XOR2_X1 \MCInst_MC1_v3_2Inst_0_U3  ( .A(\MCInst_MC1_v3_2 [3]), .B(
        \Red_MCInst_MC1_v3_3 [2]), .Z(\MCInst_MC1_v3_2 [0]) );
  XNOR2_X1 \MCInst_MC1_v3_3Inst_0_U4  ( .A(\MCInst_MC1_v3_3Inst_0_n2 ), .B(
        \Red_MCInst_MC1_v3_3 [2]), .ZN(\MCInst_MC1_v3_3 [0]) );
  XNOR2_X1 \MCInst_MC1_v3_3Inst_0_U3  ( .A(\Red_MCInst_MC1_v3_1 [2]), .B(
        \MCInst_MC1_v3_2 [3]), .ZN(\MCInst_MC1_v3_3Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC1_v0_0Inst_1_U3  ( .A(\MCInst_MC1_v0_3 [3]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\MCInst_MC1_v0_0 [1]) );
  XOR2_X1 \MCInst_MC1_v0_1Inst_1_U3  ( .A(\Red_MCInst_MC1_v0_2 [2]), .B(
        \MCInst_MC1_v0_3 [3]), .Z(\MCInst_MC1_v0_1 [1]) );
  XNOR2_X1 \MCInst_MC1_v0_2Inst_1_U4  ( .A(\MCInst_MC1_v0_2Inst_1_n2 ), .B(
        \MCInst_MC1_v0_3 [3]), .ZN(\MCInst_MC1_v0_2 [1]) );
  XNOR2_X1 \MCInst_MC1_v0_2Inst_1_U3  ( .A(\Red_MCInst_MC1_v0_1 [0]), .B(
        \Red_MCInst_MC1_v0_0 [0]), .ZN(\MCInst_MC1_v0_2Inst_1_n2 ) );
  XOR2_X1 \MCInst_MC1_v0_3Inst_1_U3  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\MCInst_MC1_v0_3 [1]) );
  XOR2_X1 \MCInst_MC1_v1_1Inst_1_U3  ( .A(\MCInst_MC1_v1_0 [0]), .B(
        \MCInst_MC1_v1_3 [3]), .Z(\MCInst_MC1_v1_1 [1]) );
  XOR2_X1 \MCInst_MC1_v1_2Inst_1_U3  ( .A(\MCInst_MC1_v1_0 [0]), .B(
        \Red_MCInst_MC1_v1_2 [1]), .Z(\MCInst_MC1_v1_2 [1]) );
  XOR2_X1 \MCInst_MC1_v1_3Inst_1_U3  ( .A(\MCInst_MC1_v1_0 [0]), .B(
        \Red_MCInst_MC1_v1_1 [2]), .Z(\MCInst_MC1_v1_3 [1]) );
  XOR2_X1 \MCInst_MC1_v2_0Inst_1_U3  ( .A(\Red_MCInst_MC1_v2_1 [1]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\MCInst_MC1_v2_0 [1]) );
  XNOR2_X1 \MCInst_MC1_v2_1Inst_1_U4  ( .A(\MCInst_MC1_v2_1Inst_1_n2 ), .B(
        \MCInst_MC1_v2_0 [3]), .ZN(\MCInst_MC1_v2_1 [1]) );
  XNOR2_X1 \MCInst_MC1_v2_1Inst_1_U3  ( .A(\Red_MCInst_MC1_v2_2 [1]), .B(
        \MCInst_MC1_v2_0 [2]), .ZN(\MCInst_MC1_v2_1Inst_1_n2 ) );
  XNOR2_X1 \MCInst_MC1_v2_2Inst_1_U5  ( .A(\MCInst_MC1_v2_2Inst_1_n4 ), .B(
        \MCInst_MC1_v2_2Inst_1_n3 ), .ZN(\MCInst_MC1_v2_2 [1]) );
  XNOR2_X1 \MCInst_MC1_v2_2Inst_1_U4  ( .A(\MCInst_MC1_v2_0 [2]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\MCInst_MC1_v2_2Inst_1_n3 ) );
  XOR2_X1 \MCInst_MC1_v2_2Inst_1_U3  ( .A(\MCInst_MC1_v2_0 [3]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\MCInst_MC1_v2_2Inst_1_n4 ) );
  XOR2_X1 \MCInst_MC1_v3_0Inst_1_U3  ( .A(\MCInst_MC1_v3_2 [3]), .B(
        \Red_MCInst_MC1_v3_1 [2]), .Z(\MCInst_MC1_v3_0 [1]) );
  XOR2_X1 \MCInst_MC1_v3_1Inst_1_U3  ( .A(\MCInst_MC1_v3_2 [3]), .B(
        \MCInst_MC1_v3_0 [3]), .Z(\MCInst_MC1_v3_1 [1]) );
  XNOR2_X1 \MCInst_MC1_v3_3Inst_1_U4  ( .A(\MCInst_MC1_v3_3Inst_1_n2 ), .B(
        \MCInst_MC1_v3_0 [3]), .ZN(\MCInst_MC1_v3_3 [1]) );
  XNOR2_X1 \MCInst_MC1_v3_3Inst_1_U3  ( .A(\Red_MCInst_MC1_v3_1 [2]), .B(
        \MCInst_MC1_v3_2 [3]), .ZN(\MCInst_MC1_v3_3Inst_1_n2 ) );
  XOR2_X1 \MCInst_MC1_v0_0Inst_2_U3  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\MCInst_MC1_v0_0 [2]) );
  XOR2_X1 \MCInst_MC1_v0_1Inst_2_U3  ( .A(\MCInst_MC1_v0_3 [3]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\MCInst_MC1_v0_1 [2]) );
  XOR2_X1 \MCInst_MC1_v0_2Inst_2_U3  ( .A(\Red_MCInst_MC1_v0_2 [2]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\MCInst_MC1_v0_2 [2]) );
  XNOR2_X1 \MCInst_MC1_v1_1Inst_2_U4  ( .A(\MCInst_MC1_v1_1Inst_2_n2 ), .B(
        \Red_MCInst_MC1_v1_2 [1]), .ZN(\MCInst_MC1_v1_1 [2]) );
  XNOR2_X1 \MCInst_MC1_v1_1Inst_2_U3  ( .A(\Red_MCInst_MC1_v1_1 [2]), .B(
        \MCInst_MC1_v1_0 [0]), .ZN(\MCInst_MC1_v1_1Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC1_v1_2Inst_2_U4  ( .A(\MCInst_MC1_v1_2Inst_2_n2 ), .B(
        \Red_MCInst_MC1_v1_2 [1]), .ZN(\MCInst_MC1_v1_2 [2]) );
  XNOR2_X1 \MCInst_MC1_v1_2Inst_2_U3  ( .A(\MCInst_MC1_v1_3 [3]), .B(
        \MCInst_MC1_v1_0 [0]), .ZN(\MCInst_MC1_v1_2Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC1_v2_1Inst_2_U4  ( .A(\MCInst_MC1_v2_1Inst_2_n2 ), .B(
        \MCInst_MC1_v2_0 [3]), .ZN(\MCInst_MC1_v2_1 [2]) );
  XNOR2_X1 \MCInst_MC1_v2_1Inst_2_U3  ( .A(\Red_MCInst_MC1_v2_2 [1]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\MCInst_MC1_v2_1Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC1_v2_2Inst_2_U4  ( .A(\MCInst_MC1_v2_2Inst_2_n2 ), .B(
        \MCInst_MC1_v2_0 [3]), .ZN(\MCInst_MC1_v2_2 [2]) );
  XNOR2_X1 \MCInst_MC1_v2_2Inst_2_U3  ( .A(\Red_MCInst_MC1_v2_2 [1]), .B(
        \MCInst_MC1_v2_0 [2]), .ZN(\MCInst_MC1_v2_2Inst_2_n2 ) );
  XOR2_X1 \MCInst_MC1_v2_3Inst_2_U3  ( .A(\Red_MCInst_MC1_v2_1 [1]), .B(
        \MCInst_MC1_v2_0 [2]), .Z(\MCInst_MC1_v2_3 [2]) );
  XNOR2_X1 \MCInst_MC1_v3_1Inst_2_U4  ( .A(\MCInst_MC1_v3_1Inst_2_n2 ), .B(
        \Red_MCInst_MC1_v3_3 [2]), .ZN(\MCInst_MC1_v3_1 [2]) );
  XNOR2_X1 \MCInst_MC1_v3_1Inst_2_U3  ( .A(\Red_MCInst_MC1_v3_1 [2]), .B(
        \MCInst_MC1_v3_2 [3]), .ZN(\MCInst_MC1_v3_1Inst_2_n2 ) );
  XOR2_X1 \MCInst_MC1_v3_3Inst_2_U3  ( .A(\Red_MCInst_MC1_v3_3 [2]), .B(
        \Red_MCInst_MC1_v3_1 [2]), .Z(\MCInst_MC1_v3_3 [2]) );
  XOR2_X1 \MCInst_MC1_v0_1Inst_3_U3  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\MCInst_MC1_v0_1 [3]) );
  XOR2_X1 \MCInst_MC1_v0_2Inst_3_U3  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(
        \MCInst_MC1_v0_3 [3]), .Z(\MCInst_MC1_v0_2 [3]) );
  XOR2_X1 \MCInst_MC1_v1_1Inst_3_U3  ( .A(\Red_MCInst_MC1_v1_2 [1]), .B(
        \MCInst_MC1_v1_3 [3]), .Z(\MCInst_MC1_v1_1 [3]) );
  XNOR2_X1 \MCInst_MC1_v1_2Inst_3_U5  ( .A(\MCInst_MC1_v1_2Inst_3_n4 ), .B(
        \MCInst_MC1_v1_2Inst_3_n3 ), .ZN(\MCInst_MC1_v1_2 [3]) );
  XNOR2_X1 \MCInst_MC1_v1_2Inst_3_U4  ( .A(\Red_MCInst_MC1_v1_2 [1]), .B(
        \MCInst_MC1_v1_0 [0]), .ZN(\MCInst_MC1_v1_2Inst_3_n3 ) );
  XOR2_X1 \MCInst_MC1_v1_2Inst_3_U3  ( .A(\MCInst_MC1_v1_3 [3]), .B(
        \Red_MCInst_MC1_v1_1 [2]), .Z(\MCInst_MC1_v1_2Inst_3_n4 ) );
  XOR2_X1 \MCInst_MC1_v2_1Inst_3_U3  ( .A(\MCInst_MC1_v2_0 [2]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\MCInst_MC1_v2_1 [3]) );
  XNOR2_X1 \MCInst_MC1_v2_2Inst_3_U4  ( .A(\MCInst_MC1_v2_2Inst_3_n2 ), .B(
        \MCInst_MC1_v2_0 [3]), .ZN(\MCInst_MC1_v2_2 [3]) );
  XNOR2_X1 \MCInst_MC1_v2_2Inst_3_U3  ( .A(\Red_MCInst_MC1_v2_2 [1]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\MCInst_MC1_v2_2Inst_3_n2 ) );
  XNOR2_X1 \MCInst_MC1_v2_3Inst_3_U4  ( .A(\MCInst_MC1_v2_3Inst_3_n2 ), .B(
        \MCInst_MC1_v2_0 [2]), .ZN(\MCInst_MC1_v2_3 [3]) );
  XNOR2_X1 \MCInst_MC1_v2_3Inst_3_U3  ( .A(\MCInst_MC1_v2_0 [3]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\MCInst_MC1_v2_3Inst_3_n2 ) );
  XOR2_X1 \MCInst_MC1_v3_1Inst_3_U3  ( .A(\Red_MCInst_MC1_v3_3 [2]), .B(
        \MCInst_MC1_v3_0 [3]), .Z(\MCInst_MC1_v3_1 [3]) );
  XOR2_X1 \MCInst_MC1_v3_3Inst_3_U3  ( .A(\MCInst_MC1_v3_2 [3]), .B(
        \MCInst_MC1_v3_0 [3]), .Z(\MCInst_MC1_v3_3 [3]) );
  XNOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC1_r0Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC1_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[56]) );
  XNOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_0_U2  ( .A(\Red_MCInst_MC1_v3_1 [2]), 
        .B(\Red_MCInst_MC1_v2_2 [1]), .ZN(\MCInst_MC1_r0Inst_XORInst_0_0_n4 )
         );
  XOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_0_U1  ( .A(\MCInst_MC1_v0_3 [3]), .B(
        \MCInst_MC1_v1_0 [0]), .Z(\MCInst_MC1_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC1_r0Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC1_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[57]) );
  XNOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_1_U2  ( .A(\MCInst_MC1_v3_0 [1]), .B(
        \MCInst_MC1_v2_0 [1]), .ZN(\MCInst_MC1_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_1_U1  ( .A(\MCInst_MC1_v0_0 [1]), .B(
        \Red_MCInst_MC1_v1_2 [1]), .Z(\MCInst_MC1_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC1_r0Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC1_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[58]) );
  XNOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_2_U2  ( .A(\Red_MCInst_MC1_v3_3 [2]), 
        .B(\MCInst_MC1_v2_0 [2]), .ZN(\MCInst_MC1_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_2_U1  ( .A(\MCInst_MC1_v0_0 [2]), .B(
        \MCInst_MC1_v1_3 [3]), .Z(\MCInst_MC1_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC1_r0Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC1_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[59]) );
  XNOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_3_U2  ( .A(\MCInst_MC1_v3_0 [3]), .B(
        \MCInst_MC1_v2_0 [3]), .ZN(\MCInst_MC1_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_3_U1  ( .A(\Red_MCInst_MC1_v0_2 [2]), 
        .B(\Red_MCInst_MC1_v1_1 [2]), .Z(\MCInst_MC1_r0Inst_XORInst_0_3_n5 )
         );
  XNOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC1_r1Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC1_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[40]) );
  XNOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_0_U2  ( .A(\MCInst_MC1_v3_1 [0]), .B(
        \MCInst_MC1_v2_1 [0]), .ZN(\MCInst_MC1_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC1_v0_2 [2]), 
        .B(\MCInst_MC1_v1_1 [0]), .Z(\MCInst_MC1_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC1_r1Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC1_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[41]) );
  XNOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_1_U2  ( .A(\MCInst_MC1_v3_1 [1]), .B(
        \MCInst_MC1_v2_1 [1]), .ZN(\MCInst_MC1_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_1_U1  ( .A(\MCInst_MC1_v0_1 [1]), .B(
        \MCInst_MC1_v1_1 [1]), .Z(\MCInst_MC1_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC1_r1Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC1_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[42]) );
  XNOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_2_U2  ( .A(\MCInst_MC1_v3_1 [2]), .B(
        \MCInst_MC1_v2_1 [2]), .ZN(\MCInst_MC1_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_2_U1  ( .A(\MCInst_MC1_v0_1 [2]), .B(
        \MCInst_MC1_v1_1 [2]), .Z(\MCInst_MC1_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC1_r1Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC1_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[43]) );
  XNOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_3_U2  ( .A(\MCInst_MC1_v3_1 [3]), .B(
        \MCInst_MC1_v2_1 [3]), .ZN(\MCInst_MC1_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_3_U1  ( .A(\MCInst_MC1_v0_1 [3]), .B(
        \MCInst_MC1_v1_1 [3]), .Z(\MCInst_MC1_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC1_r2Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC1_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[24]) );
  XNOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_0_U2  ( .A(\MCInst_MC1_v3_2 [0]), .B(
        \MCInst_MC1_v2_2 [0]), .ZN(\MCInst_MC1_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_0_U1  ( .A(\MCInst_MC1_v0_2 [0]), .B(
        \MCInst_MC1_v1_2 [0]), .Z(\MCInst_MC1_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC1_r2Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC1_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[25]) );
  XNOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_1_U2  ( .A(\MCInst_MC1_v3_0 [3]), .B(
        \MCInst_MC1_v2_2 [1]), .ZN(\MCInst_MC1_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_1_U1  ( .A(\MCInst_MC1_v0_2 [1]), .B(
        \MCInst_MC1_v1_2 [1]), .Z(\MCInst_MC1_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC1_r2Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC1_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[26]) );
  XNOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_2_U2  ( .A(\Red_MCInst_MC1_v3_1 [2]), 
        .B(\MCInst_MC1_v2_2 [2]), .ZN(\MCInst_MC1_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_2_U1  ( .A(\MCInst_MC1_v0_2 [2]), .B(
        \MCInst_MC1_v1_2 [2]), .Z(\MCInst_MC1_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC1_r2Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC1_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[27]) );
  XNOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_3_U2  ( .A(\MCInst_MC1_v3_2 [3]), .B(
        \MCInst_MC1_v2_2 [3]), .ZN(\MCInst_MC1_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_3_U1  ( .A(\MCInst_MC1_v0_2 [3]), .B(
        \MCInst_MC1_v1_2 [3]), .Z(\MCInst_MC1_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC1_r3Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC1_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[8]) );
  XNOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_0_U2  ( .A(\MCInst_MC1_v3_3 [0]), .B(
        \MCInst_MC1_v2_3 [0]), .ZN(\MCInst_MC1_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC1_v0_1 [0]), 
        .B(\Red_MCInst_MC1_v1_1 [2]), .Z(\MCInst_MC1_r3Inst_XORInst_0_0_n5 )
         );
  XNOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC1_r3Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC1_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[9]) );
  XNOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_1_U2  ( .A(\MCInst_MC1_v3_3 [1]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\MCInst_MC1_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_1_U1  ( .A(\MCInst_MC1_v0_3 [1]), .B(
        \MCInst_MC1_v1_3 [1]), .Z(\MCInst_MC1_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC1_r3Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC1_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[10]) );
  XNOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_2_U2  ( .A(\MCInst_MC1_v3_3 [2]), .B(
        \MCInst_MC1_v2_3 [2]), .ZN(\MCInst_MC1_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC1_v0_2 [2]), 
        .B(\Red_MCInst_MC1_v1_2 [1]), .Z(\MCInst_MC1_r3Inst_XORInst_0_2_n5 )
         );
  XNOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC1_r3Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC1_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[11]) );
  XNOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_3_U2  ( .A(\MCInst_MC1_v3_3 [3]), .B(
        \MCInst_MC1_v2_3 [3]), .ZN(\MCInst_MC1_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_3_U1  ( .A(\MCInst_MC1_v0_3 [3]), .B(
        \MCInst_MC1_v1_3 [3]), .Z(\MCInst_MC1_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC2_v0_2Inst_0_U4  ( .A(\MCInst_MC2_v0_2Inst_0_n2 ), .B(
        \Red_MCInst_MC2_v0_2 [2]), .ZN(\MCInst_MC2_v0_2 [0]) );
  XNOR2_X1 \MCInst_MC2_v0_2Inst_0_U3  ( .A(\Red_MCInst_MC2_v0_1 [0]), .B(
        \Red_MCInst_MC2_v0_0 [0]), .ZN(\MCInst_MC2_v0_2Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC2_v1_1Inst_0_U3  ( .A(\MCInst_MC2_v1_3 [3]), .B(
        \Red_MCInst_MC2_v1_1 [2]), .Z(\MCInst_MC2_v1_1 [0]) );
  XNOR2_X1 \MCInst_MC2_v1_2Inst_0_U4  ( .A(\MCInst_MC2_v1_2Inst_0_n2 ), .B(
        \MCInst_MC2_v1_3 [3]), .ZN(\MCInst_MC2_v1_2 [0]) );
  XNOR2_X1 \MCInst_MC2_v1_2Inst_0_U3  ( .A(\Red_MCInst_MC2_v1_1 [2]), .B(
        \Red_MCInst_MC2_v1_2 [1]), .ZN(\MCInst_MC2_v1_2Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC2_v2_1Inst_0_U3  ( .A(\Red_MCInst_MC2_v2_1 [1]), .B(
        \MCInst_MC2_v2_0 [3]), .Z(\MCInst_MC2_v2_1 [0]) );
  XOR2_X1 \MCInst_MC2_v2_2Inst_0_U3  ( .A(\MCInst_MC2_v2_0 [2]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\MCInst_MC2_v2_2 [0]) );
  XNOR2_X1 \MCInst_MC2_v2_3Inst_0_U5  ( .A(\MCInst_MC2_v2_3Inst_0_n4 ), .B(
        \MCInst_MC2_v2_3Inst_0_n3 ), .ZN(\MCInst_MC2_v2_3 [0]) );
  XNOR2_X1 \MCInst_MC2_v2_3Inst_0_U4  ( .A(\MCInst_MC2_v2_0 [2]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\MCInst_MC2_v2_3Inst_0_n3 ) );
  XOR2_X1 \MCInst_MC2_v2_3Inst_0_U3  ( .A(\MCInst_MC2_v2_0 [3]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\MCInst_MC2_v2_3Inst_0_n4 ) );
  XOR2_X1 \MCInst_MC2_v3_1Inst_0_U3  ( .A(\MCInst_MC2_v3_0 [3]), .B(
        \Red_MCInst_MC2_v3_1 [2]), .Z(\MCInst_MC2_v3_1 [0]) );
  XOR2_X1 \MCInst_MC2_v3_2Inst_0_U3  ( .A(\MCInst_MC2_v3_2 [3]), .B(
        \Red_MCInst_MC2_v3_3 [2]), .Z(\MCInst_MC2_v3_2 [0]) );
  XNOR2_X1 \MCInst_MC2_v3_3Inst_0_U4  ( .A(\MCInst_MC2_v3_3Inst_0_n2 ), .B(
        \Red_MCInst_MC2_v3_3 [2]), .ZN(\MCInst_MC2_v3_3 [0]) );
  XNOR2_X1 \MCInst_MC2_v3_3Inst_0_U3  ( .A(\Red_MCInst_MC2_v3_1 [2]), .B(
        \MCInst_MC2_v3_2 [3]), .ZN(\MCInst_MC2_v3_3Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC2_v0_0Inst_1_U3  ( .A(\MCInst_MC2_v0_3 [3]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\MCInst_MC2_v0_0 [1]) );
  XOR2_X1 \MCInst_MC2_v0_1Inst_1_U3  ( .A(\Red_MCInst_MC2_v0_2 [2]), .B(
        \MCInst_MC2_v0_3 [3]), .Z(\MCInst_MC2_v0_1 [1]) );
  XNOR2_X1 \MCInst_MC2_v0_2Inst_1_U4  ( .A(\MCInst_MC2_v0_2Inst_1_n2 ), .B(
        \MCInst_MC2_v0_3 [3]), .ZN(\MCInst_MC2_v0_2 [1]) );
  XNOR2_X1 \MCInst_MC2_v0_2Inst_1_U3  ( .A(\Red_MCInst_MC2_v0_1 [0]), .B(
        \Red_MCInst_MC2_v0_0 [0]), .ZN(\MCInst_MC2_v0_2Inst_1_n2 ) );
  XOR2_X1 \MCInst_MC2_v0_3Inst_1_U3  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\MCInst_MC2_v0_3 [1]) );
  XOR2_X1 \MCInst_MC2_v1_1Inst_1_U3  ( .A(\MCInst_MC2_v1_0 [0]), .B(
        \MCInst_MC2_v1_3 [3]), .Z(\MCInst_MC2_v1_1 [1]) );
  XOR2_X1 \MCInst_MC2_v1_2Inst_1_U3  ( .A(\MCInst_MC2_v1_0 [0]), .B(
        \Red_MCInst_MC2_v1_2 [1]), .Z(\MCInst_MC2_v1_2 [1]) );
  XOR2_X1 \MCInst_MC2_v1_3Inst_1_U3  ( .A(\MCInst_MC2_v1_0 [0]), .B(
        \Red_MCInst_MC2_v1_1 [2]), .Z(\MCInst_MC2_v1_3 [1]) );
  XOR2_X1 \MCInst_MC2_v2_0Inst_1_U3  ( .A(\Red_MCInst_MC2_v2_1 [1]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\MCInst_MC2_v2_0 [1]) );
  XNOR2_X1 \MCInst_MC2_v2_1Inst_1_U4  ( .A(\MCInst_MC2_v2_1Inst_1_n2 ), .B(
        \MCInst_MC2_v2_0 [3]), .ZN(\MCInst_MC2_v2_1 [1]) );
  XNOR2_X1 \MCInst_MC2_v2_1Inst_1_U3  ( .A(\Red_MCInst_MC2_v2_2 [1]), .B(
        \MCInst_MC2_v2_0 [2]), .ZN(\MCInst_MC2_v2_1Inst_1_n2 ) );
  XNOR2_X1 \MCInst_MC2_v2_2Inst_1_U5  ( .A(\MCInst_MC2_v2_2Inst_1_n4 ), .B(
        \MCInst_MC2_v2_2Inst_1_n3 ), .ZN(\MCInst_MC2_v2_2 [1]) );
  XNOR2_X1 \MCInst_MC2_v2_2Inst_1_U4  ( .A(\MCInst_MC2_v2_0 [2]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\MCInst_MC2_v2_2Inst_1_n3 ) );
  XOR2_X1 \MCInst_MC2_v2_2Inst_1_U3  ( .A(\MCInst_MC2_v2_0 [3]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\MCInst_MC2_v2_2Inst_1_n4 ) );
  XOR2_X1 \MCInst_MC2_v3_0Inst_1_U3  ( .A(\MCInst_MC2_v3_2 [3]), .B(
        \Red_MCInst_MC2_v3_1 [2]), .Z(\MCInst_MC2_v3_0 [1]) );
  XOR2_X1 \MCInst_MC2_v3_1Inst_1_U3  ( .A(\MCInst_MC2_v3_2 [3]), .B(
        \MCInst_MC2_v3_0 [3]), .Z(\MCInst_MC2_v3_1 [1]) );
  XNOR2_X1 \MCInst_MC2_v3_3Inst_1_U4  ( .A(\MCInst_MC2_v3_3Inst_1_n2 ), .B(
        \MCInst_MC2_v3_0 [3]), .ZN(\MCInst_MC2_v3_3 [1]) );
  XNOR2_X1 \MCInst_MC2_v3_3Inst_1_U3  ( .A(\Red_MCInst_MC2_v3_1 [2]), .B(
        \MCInst_MC2_v3_2 [3]), .ZN(\MCInst_MC2_v3_3Inst_1_n2 ) );
  XOR2_X1 \MCInst_MC2_v0_0Inst_2_U3  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\MCInst_MC2_v0_0 [2]) );
  XOR2_X1 \MCInst_MC2_v0_1Inst_2_U3  ( .A(\MCInst_MC2_v0_3 [3]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\MCInst_MC2_v0_1 [2]) );
  XOR2_X1 \MCInst_MC2_v0_2Inst_2_U3  ( .A(\Red_MCInst_MC2_v0_2 [2]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\MCInst_MC2_v0_2 [2]) );
  XNOR2_X1 \MCInst_MC2_v1_1Inst_2_U4  ( .A(\MCInst_MC2_v1_1Inst_2_n2 ), .B(
        \Red_MCInst_MC2_v1_2 [1]), .ZN(\MCInst_MC2_v1_1 [2]) );
  XNOR2_X1 \MCInst_MC2_v1_1Inst_2_U3  ( .A(\Red_MCInst_MC2_v1_1 [2]), .B(
        \MCInst_MC2_v1_0 [0]), .ZN(\MCInst_MC2_v1_1Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC2_v1_2Inst_2_U4  ( .A(\MCInst_MC2_v1_2Inst_2_n2 ), .B(
        \Red_MCInst_MC2_v1_2 [1]), .ZN(\MCInst_MC2_v1_2 [2]) );
  XNOR2_X1 \MCInst_MC2_v1_2Inst_2_U3  ( .A(\MCInst_MC2_v1_3 [3]), .B(
        \MCInst_MC2_v1_0 [0]), .ZN(\MCInst_MC2_v1_2Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC2_v2_1Inst_2_U4  ( .A(\MCInst_MC2_v2_1Inst_2_n2 ), .B(
        \MCInst_MC2_v2_0 [3]), .ZN(\MCInst_MC2_v2_1 [2]) );
  XNOR2_X1 \MCInst_MC2_v2_1Inst_2_U3  ( .A(\Red_MCInst_MC2_v2_2 [1]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\MCInst_MC2_v2_1Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC2_v2_2Inst_2_U4  ( .A(\MCInst_MC2_v2_2Inst_2_n2 ), .B(
        \MCInst_MC2_v2_0 [3]), .ZN(\MCInst_MC2_v2_2 [2]) );
  XNOR2_X1 \MCInst_MC2_v2_2Inst_2_U3  ( .A(\Red_MCInst_MC2_v2_2 [1]), .B(
        \MCInst_MC2_v2_0 [2]), .ZN(\MCInst_MC2_v2_2Inst_2_n2 ) );
  XOR2_X1 \MCInst_MC2_v2_3Inst_2_U3  ( .A(\Red_MCInst_MC2_v2_1 [1]), .B(
        \MCInst_MC2_v2_0 [2]), .Z(\MCInst_MC2_v2_3 [2]) );
  XNOR2_X1 \MCInst_MC2_v3_1Inst_2_U4  ( .A(\MCInst_MC2_v3_1Inst_2_n2 ), .B(
        \Red_MCInst_MC2_v3_3 [2]), .ZN(\MCInst_MC2_v3_1 [2]) );
  XNOR2_X1 \MCInst_MC2_v3_1Inst_2_U3  ( .A(\Red_MCInst_MC2_v3_1 [2]), .B(
        \MCInst_MC2_v3_2 [3]), .ZN(\MCInst_MC2_v3_1Inst_2_n2 ) );
  XOR2_X1 \MCInst_MC2_v3_3Inst_2_U3  ( .A(\Red_MCInst_MC2_v3_3 [2]), .B(
        \Red_MCInst_MC2_v3_1 [2]), .Z(\MCInst_MC2_v3_3 [2]) );
  XOR2_X1 \MCInst_MC2_v0_1Inst_3_U3  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\MCInst_MC2_v0_1 [3]) );
  XOR2_X1 \MCInst_MC2_v0_2Inst_3_U3  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(
        \MCInst_MC2_v0_3 [3]), .Z(\MCInst_MC2_v0_2 [3]) );
  XOR2_X1 \MCInst_MC2_v1_1Inst_3_U3  ( .A(\Red_MCInst_MC2_v1_2 [1]), .B(
        \MCInst_MC2_v1_3 [3]), .Z(\MCInst_MC2_v1_1 [3]) );
  XNOR2_X1 \MCInst_MC2_v1_2Inst_3_U5  ( .A(\MCInst_MC2_v1_2Inst_3_n4 ), .B(
        \MCInst_MC2_v1_2Inst_3_n3 ), .ZN(\MCInst_MC2_v1_2 [3]) );
  XNOR2_X1 \MCInst_MC2_v1_2Inst_3_U4  ( .A(\Red_MCInst_MC2_v1_2 [1]), .B(
        \MCInst_MC2_v1_0 [0]), .ZN(\MCInst_MC2_v1_2Inst_3_n3 ) );
  XOR2_X1 \MCInst_MC2_v1_2Inst_3_U3  ( .A(\MCInst_MC2_v1_3 [3]), .B(
        \Red_MCInst_MC2_v1_1 [2]), .Z(\MCInst_MC2_v1_2Inst_3_n4 ) );
  XOR2_X1 \MCInst_MC2_v2_1Inst_3_U3  ( .A(\MCInst_MC2_v2_0 [2]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\MCInst_MC2_v2_1 [3]) );
  XNOR2_X1 \MCInst_MC2_v2_2Inst_3_U4  ( .A(\MCInst_MC2_v2_2Inst_3_n2 ), .B(
        \MCInst_MC2_v2_0 [3]), .ZN(\MCInst_MC2_v2_2 [3]) );
  XNOR2_X1 \MCInst_MC2_v2_2Inst_3_U3  ( .A(\Red_MCInst_MC2_v2_2 [1]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\MCInst_MC2_v2_2Inst_3_n2 ) );
  XNOR2_X1 \MCInst_MC2_v2_3Inst_3_U4  ( .A(\MCInst_MC2_v2_3Inst_3_n2 ), .B(
        \MCInst_MC2_v2_0 [2]), .ZN(\MCInst_MC2_v2_3 [3]) );
  XNOR2_X1 \MCInst_MC2_v2_3Inst_3_U3  ( .A(\MCInst_MC2_v2_0 [3]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\MCInst_MC2_v2_3Inst_3_n2 ) );
  XOR2_X1 \MCInst_MC2_v3_1Inst_3_U3  ( .A(\Red_MCInst_MC2_v3_3 [2]), .B(
        \MCInst_MC2_v3_0 [3]), .Z(\MCInst_MC2_v3_1 [3]) );
  XOR2_X1 \MCInst_MC2_v3_3Inst_3_U3  ( .A(\MCInst_MC2_v3_2 [3]), .B(
        \MCInst_MC2_v3_0 [3]), .Z(\MCInst_MC2_v3_3 [3]) );
  XNOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC2_r0Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC2_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[52]) );
  XNOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_0_U2  ( .A(\Red_MCInst_MC2_v3_1 [2]), 
        .B(\Red_MCInst_MC2_v2_2 [1]), .ZN(\MCInst_MC2_r0Inst_XORInst_0_0_n4 )
         );
  XOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_0_U1  ( .A(\MCInst_MC2_v0_3 [3]), .B(
        \MCInst_MC2_v1_0 [0]), .Z(\MCInst_MC2_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC2_r0Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC2_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[53]) );
  XNOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_1_U2  ( .A(\MCInst_MC2_v3_0 [1]), .B(
        \MCInst_MC2_v2_0 [1]), .ZN(\MCInst_MC2_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_1_U1  ( .A(\MCInst_MC2_v0_0 [1]), .B(
        \Red_MCInst_MC2_v1_2 [1]), .Z(\MCInst_MC2_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC2_r0Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC2_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[54]) );
  XNOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_2_U2  ( .A(\Red_MCInst_MC2_v3_3 [2]), 
        .B(\MCInst_MC2_v2_0 [2]), .ZN(\MCInst_MC2_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_2_U1  ( .A(\MCInst_MC2_v0_0 [2]), .B(
        \MCInst_MC2_v1_3 [3]), .Z(\MCInst_MC2_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC2_r0Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC2_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[55]) );
  XNOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_3_U2  ( .A(\MCInst_MC2_v3_0 [3]), .B(
        \MCInst_MC2_v2_0 [3]), .ZN(\MCInst_MC2_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_3_U1  ( .A(\Red_MCInst_MC2_v0_2 [2]), 
        .B(\Red_MCInst_MC2_v1_1 [2]), .Z(\MCInst_MC2_r0Inst_XORInst_0_3_n5 )
         );
  XNOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC2_r1Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC2_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[36]) );
  XNOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_0_U2  ( .A(\MCInst_MC2_v3_1 [0]), .B(
        \MCInst_MC2_v2_1 [0]), .ZN(\MCInst_MC2_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC2_v0_2 [2]), 
        .B(\MCInst_MC2_v1_1 [0]), .Z(\MCInst_MC2_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC2_r1Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC2_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[37]) );
  XNOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_1_U2  ( .A(\MCInst_MC2_v3_1 [1]), .B(
        \MCInst_MC2_v2_1 [1]), .ZN(\MCInst_MC2_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_1_U1  ( .A(\MCInst_MC2_v0_1 [1]), .B(
        \MCInst_MC2_v1_1 [1]), .Z(\MCInst_MC2_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC2_r1Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC2_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[38]) );
  XNOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_2_U2  ( .A(\MCInst_MC2_v3_1 [2]), .B(
        \MCInst_MC2_v2_1 [2]), .ZN(\MCInst_MC2_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_2_U1  ( .A(\MCInst_MC2_v0_1 [2]), .B(
        \MCInst_MC2_v1_1 [2]), .Z(\MCInst_MC2_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC2_r1Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC2_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[39]) );
  XNOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_3_U2  ( .A(\MCInst_MC2_v3_1 [3]), .B(
        \MCInst_MC2_v2_1 [3]), .ZN(\MCInst_MC2_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_3_U1  ( .A(\MCInst_MC2_v0_1 [3]), .B(
        \MCInst_MC2_v1_1 [3]), .Z(\MCInst_MC2_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC2_r2Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC2_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[20]) );
  XNOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_0_U2  ( .A(\MCInst_MC2_v3_2 [0]), .B(
        \MCInst_MC2_v2_2 [0]), .ZN(\MCInst_MC2_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_0_U1  ( .A(\MCInst_MC2_v0_2 [0]), .B(
        \MCInst_MC2_v1_2 [0]), .Z(\MCInst_MC2_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC2_r2Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC2_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[21]) );
  XNOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_1_U2  ( .A(\MCInst_MC2_v3_0 [3]), .B(
        \MCInst_MC2_v2_2 [1]), .ZN(\MCInst_MC2_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_1_U1  ( .A(\MCInst_MC2_v0_2 [1]), .B(
        \MCInst_MC2_v1_2 [1]), .Z(\MCInst_MC2_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC2_r2Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC2_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[22]) );
  XNOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_2_U2  ( .A(\Red_MCInst_MC2_v3_1 [2]), 
        .B(\MCInst_MC2_v2_2 [2]), .ZN(\MCInst_MC2_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_2_U1  ( .A(\MCInst_MC2_v0_2 [2]), .B(
        \MCInst_MC2_v1_2 [2]), .Z(\MCInst_MC2_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC2_r2Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC2_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[23]) );
  XNOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_3_U2  ( .A(\MCInst_MC2_v3_2 [3]), .B(
        \MCInst_MC2_v2_2 [3]), .ZN(\MCInst_MC2_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_3_U1  ( .A(\MCInst_MC2_v0_2 [3]), .B(
        \MCInst_MC2_v1_2 [3]), .Z(\MCInst_MC2_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC2_r3Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC2_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[4]) );
  XNOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_0_U2  ( .A(\MCInst_MC2_v3_3 [0]), .B(
        \MCInst_MC2_v2_3 [0]), .ZN(\MCInst_MC2_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC2_v0_1 [0]), 
        .B(\Red_MCInst_MC2_v1_1 [2]), .Z(\MCInst_MC2_r3Inst_XORInst_0_0_n5 )
         );
  XNOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC2_r3Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC2_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[5]) );
  XNOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_1_U2  ( .A(\MCInst_MC2_v3_3 [1]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\MCInst_MC2_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_1_U1  ( .A(\MCInst_MC2_v0_3 [1]), .B(
        \MCInst_MC2_v1_3 [1]), .Z(\MCInst_MC2_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC2_r3Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC2_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[6]) );
  XNOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_2_U2  ( .A(\MCInst_MC2_v3_3 [2]), .B(
        \MCInst_MC2_v2_3 [2]), .ZN(\MCInst_MC2_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC2_v0_2 [2]), 
        .B(\Red_MCInst_MC2_v1_2 [1]), .Z(\MCInst_MC2_r3Inst_XORInst_0_2_n5 )
         );
  XNOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC2_r3Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC2_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[7]) );
  XNOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_3_U2  ( .A(\MCInst_MC2_v3_3 [3]), .B(
        \MCInst_MC2_v2_3 [3]), .ZN(\MCInst_MC2_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_3_U1  ( .A(\MCInst_MC2_v0_3 [3]), .B(
        \MCInst_MC2_v1_3 [3]), .Z(\MCInst_MC2_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC3_v0_2Inst_0_U4  ( .A(\MCInst_MC3_v0_2Inst_0_n2 ), .B(
        \Red_MCInst_MC3_v0_2 [2]), .ZN(\MCInst_MC3_v0_2 [0]) );
  XNOR2_X1 \MCInst_MC3_v0_2Inst_0_U3  ( .A(\Red_MCInst_MC3_v0_1 [0]), .B(
        \Red_MCInst_MC3_v0_0 [0]), .ZN(\MCInst_MC3_v0_2Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC3_v1_1Inst_0_U3  ( .A(\MCInst_MC3_v1_3 [3]), .B(
        \Red_MCInst_MC3_v1_1 [2]), .Z(\MCInst_MC3_v1_1 [0]) );
  XNOR2_X1 \MCInst_MC3_v1_2Inst_0_U4  ( .A(\MCInst_MC3_v1_2Inst_0_n2 ), .B(
        \MCInst_MC3_v1_3 [3]), .ZN(\MCInst_MC3_v1_2 [0]) );
  XNOR2_X1 \MCInst_MC3_v1_2Inst_0_U3  ( .A(\Red_MCInst_MC3_v1_1 [2]), .B(
        \Red_MCInst_MC3_v1_2 [1]), .ZN(\MCInst_MC3_v1_2Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC3_v2_1Inst_0_U3  ( .A(\Red_MCInst_MC3_v2_1 [1]), .B(
        \MCInst_MC3_v2_0 [3]), .Z(\MCInst_MC3_v2_1 [0]) );
  XOR2_X1 \MCInst_MC3_v2_2Inst_0_U3  ( .A(\MCInst_MC3_v2_0 [2]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\MCInst_MC3_v2_2 [0]) );
  XNOR2_X1 \MCInst_MC3_v2_3Inst_0_U5  ( .A(\MCInst_MC3_v2_3Inst_0_n4 ), .B(
        \MCInst_MC3_v2_3Inst_0_n3 ), .ZN(\MCInst_MC3_v2_3 [0]) );
  XNOR2_X1 \MCInst_MC3_v2_3Inst_0_U4  ( .A(\MCInst_MC3_v2_0 [2]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\MCInst_MC3_v2_3Inst_0_n3 ) );
  XOR2_X1 \MCInst_MC3_v2_3Inst_0_U3  ( .A(\MCInst_MC3_v2_0 [3]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\MCInst_MC3_v2_3Inst_0_n4 ) );
  XOR2_X1 \MCInst_MC3_v3_1Inst_0_U3  ( .A(\MCInst_MC3_v3_0 [3]), .B(
        \Red_MCInst_MC3_v3_1 [2]), .Z(\MCInst_MC3_v3_1 [0]) );
  XOR2_X1 \MCInst_MC3_v3_2Inst_0_U3  ( .A(\MCInst_MC3_v3_2 [3]), .B(
        \Red_MCInst_MC3_v3_3 [2]), .Z(\MCInst_MC3_v3_2 [0]) );
  XNOR2_X1 \MCInst_MC3_v3_3Inst_0_U4  ( .A(\MCInst_MC3_v3_3Inst_0_n2 ), .B(
        \Red_MCInst_MC3_v3_3 [2]), .ZN(\MCInst_MC3_v3_3 [0]) );
  XNOR2_X1 \MCInst_MC3_v3_3Inst_0_U3  ( .A(\Red_MCInst_MC3_v3_1 [2]), .B(
        \MCInst_MC3_v3_2 [3]), .ZN(\MCInst_MC3_v3_3Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC3_v0_0Inst_1_U3  ( .A(\MCInst_MC3_v0_3 [3]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\MCInst_MC3_v0_0 [1]) );
  XOR2_X1 \MCInst_MC3_v0_1Inst_1_U3  ( .A(\Red_MCInst_MC3_v0_2 [2]), .B(
        \MCInst_MC3_v0_3 [3]), .Z(\MCInst_MC3_v0_1 [1]) );
  XNOR2_X1 \MCInst_MC3_v0_2Inst_1_U4  ( .A(\MCInst_MC3_v0_2Inst_1_n2 ), .B(
        \MCInst_MC3_v0_3 [3]), .ZN(\MCInst_MC3_v0_2 [1]) );
  XNOR2_X1 \MCInst_MC3_v0_2Inst_1_U3  ( .A(\Red_MCInst_MC3_v0_1 [0]), .B(
        \Red_MCInst_MC3_v0_0 [0]), .ZN(\MCInst_MC3_v0_2Inst_1_n2 ) );
  XOR2_X1 \MCInst_MC3_v0_3Inst_1_U3  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\MCInst_MC3_v0_3 [1]) );
  XOR2_X1 \MCInst_MC3_v1_1Inst_1_U3  ( .A(\MCInst_MC3_v1_0 [0]), .B(
        \MCInst_MC3_v1_3 [3]), .Z(\MCInst_MC3_v1_1 [1]) );
  XOR2_X1 \MCInst_MC3_v1_2Inst_1_U3  ( .A(\MCInst_MC3_v1_0 [0]), .B(
        \Red_MCInst_MC3_v1_2 [1]), .Z(\MCInst_MC3_v1_2 [1]) );
  XOR2_X1 \MCInst_MC3_v1_3Inst_1_U3  ( .A(\MCInst_MC3_v1_0 [0]), .B(
        \Red_MCInst_MC3_v1_1 [2]), .Z(\MCInst_MC3_v1_3 [1]) );
  XOR2_X1 \MCInst_MC3_v2_0Inst_1_U3  ( .A(\Red_MCInst_MC3_v2_1 [1]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\MCInst_MC3_v2_0 [1]) );
  XNOR2_X1 \MCInst_MC3_v2_1Inst_1_U4  ( .A(\MCInst_MC3_v2_1Inst_1_n2 ), .B(
        \MCInst_MC3_v2_0 [3]), .ZN(\MCInst_MC3_v2_1 [1]) );
  XNOR2_X1 \MCInst_MC3_v2_1Inst_1_U3  ( .A(\Red_MCInst_MC3_v2_2 [1]), .B(
        \MCInst_MC3_v2_0 [2]), .ZN(\MCInst_MC3_v2_1Inst_1_n2 ) );
  XNOR2_X1 \MCInst_MC3_v2_2Inst_1_U5  ( .A(\MCInst_MC3_v2_2Inst_1_n4 ), .B(
        \MCInst_MC3_v2_2Inst_1_n3 ), .ZN(\MCInst_MC3_v2_2 [1]) );
  XNOR2_X1 \MCInst_MC3_v2_2Inst_1_U4  ( .A(\MCInst_MC3_v2_0 [2]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\MCInst_MC3_v2_2Inst_1_n3 ) );
  XOR2_X1 \MCInst_MC3_v2_2Inst_1_U3  ( .A(\MCInst_MC3_v2_0 [3]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\MCInst_MC3_v2_2Inst_1_n4 ) );
  XOR2_X1 \MCInst_MC3_v3_0Inst_1_U3  ( .A(\MCInst_MC3_v3_2 [3]), .B(
        \Red_MCInst_MC3_v3_1 [2]), .Z(\MCInst_MC3_v3_0 [1]) );
  XOR2_X1 \MCInst_MC3_v3_1Inst_1_U3  ( .A(\MCInst_MC3_v3_2 [3]), .B(
        \MCInst_MC3_v3_0 [3]), .Z(\MCInst_MC3_v3_1 [1]) );
  XNOR2_X1 \MCInst_MC3_v3_3Inst_1_U4  ( .A(\MCInst_MC3_v3_3Inst_1_n2 ), .B(
        \MCInst_MC3_v3_0 [3]), .ZN(\MCInst_MC3_v3_3 [1]) );
  XNOR2_X1 \MCInst_MC3_v3_3Inst_1_U3  ( .A(\Red_MCInst_MC3_v3_1 [2]), .B(
        \MCInst_MC3_v3_2 [3]), .ZN(\MCInst_MC3_v3_3Inst_1_n2 ) );
  XOR2_X1 \MCInst_MC3_v0_0Inst_2_U3  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\MCInst_MC3_v0_0 [2]) );
  XOR2_X1 \MCInst_MC3_v0_1Inst_2_U3  ( .A(\MCInst_MC3_v0_3 [3]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\MCInst_MC3_v0_1 [2]) );
  XOR2_X1 \MCInst_MC3_v0_2Inst_2_U3  ( .A(\Red_MCInst_MC3_v0_2 [2]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\MCInst_MC3_v0_2 [2]) );
  XNOR2_X1 \MCInst_MC3_v1_1Inst_2_U4  ( .A(\MCInst_MC3_v1_1Inst_2_n2 ), .B(
        \Red_MCInst_MC3_v1_2 [1]), .ZN(\MCInst_MC3_v1_1 [2]) );
  XNOR2_X1 \MCInst_MC3_v1_1Inst_2_U3  ( .A(\Red_MCInst_MC3_v1_1 [2]), .B(
        \MCInst_MC3_v1_0 [0]), .ZN(\MCInst_MC3_v1_1Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC3_v1_2Inst_2_U4  ( .A(\MCInst_MC3_v1_2Inst_2_n2 ), .B(
        \Red_MCInst_MC3_v1_2 [1]), .ZN(\MCInst_MC3_v1_2 [2]) );
  XNOR2_X1 \MCInst_MC3_v1_2Inst_2_U3  ( .A(\MCInst_MC3_v1_3 [3]), .B(
        \MCInst_MC3_v1_0 [0]), .ZN(\MCInst_MC3_v1_2Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC3_v2_1Inst_2_U4  ( .A(\MCInst_MC3_v2_1Inst_2_n2 ), .B(
        \MCInst_MC3_v2_0 [3]), .ZN(\MCInst_MC3_v2_1 [2]) );
  XNOR2_X1 \MCInst_MC3_v2_1Inst_2_U3  ( .A(\Red_MCInst_MC3_v2_2 [1]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\MCInst_MC3_v2_1Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC3_v2_2Inst_2_U4  ( .A(\MCInst_MC3_v2_2Inst_2_n2 ), .B(
        \MCInst_MC3_v2_0 [3]), .ZN(\MCInst_MC3_v2_2 [2]) );
  XNOR2_X1 \MCInst_MC3_v2_2Inst_2_U3  ( .A(\Red_MCInst_MC3_v2_2 [1]), .B(
        \MCInst_MC3_v2_0 [2]), .ZN(\MCInst_MC3_v2_2Inst_2_n2 ) );
  XOR2_X1 \MCInst_MC3_v2_3Inst_2_U3  ( .A(\Red_MCInst_MC3_v2_1 [1]), .B(
        \MCInst_MC3_v2_0 [2]), .Z(\MCInst_MC3_v2_3 [2]) );
  XNOR2_X1 \MCInst_MC3_v3_1Inst_2_U4  ( .A(\MCInst_MC3_v3_1Inst_2_n2 ), .B(
        \Red_MCInst_MC3_v3_3 [2]), .ZN(\MCInst_MC3_v3_1 [2]) );
  XNOR2_X1 \MCInst_MC3_v3_1Inst_2_U3  ( .A(\Red_MCInst_MC3_v3_1 [2]), .B(
        \MCInst_MC3_v3_2 [3]), .ZN(\MCInst_MC3_v3_1Inst_2_n2 ) );
  XOR2_X1 \MCInst_MC3_v3_3Inst_2_U3  ( .A(\Red_MCInst_MC3_v3_3 [2]), .B(
        \Red_MCInst_MC3_v3_1 [2]), .Z(\MCInst_MC3_v3_3 [2]) );
  XOR2_X1 \MCInst_MC3_v0_1Inst_3_U3  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\MCInst_MC3_v0_1 [3]) );
  XOR2_X1 \MCInst_MC3_v0_2Inst_3_U3  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(
        \MCInst_MC3_v0_3 [3]), .Z(\MCInst_MC3_v0_2 [3]) );
  XOR2_X1 \MCInst_MC3_v1_1Inst_3_U3  ( .A(\Red_MCInst_MC3_v1_2 [1]), .B(
        \MCInst_MC3_v1_3 [3]), .Z(\MCInst_MC3_v1_1 [3]) );
  XNOR2_X1 \MCInst_MC3_v1_2Inst_3_U5  ( .A(\MCInst_MC3_v1_2Inst_3_n4 ), .B(
        \MCInst_MC3_v1_2Inst_3_n3 ), .ZN(\MCInst_MC3_v1_2 [3]) );
  XNOR2_X1 \MCInst_MC3_v1_2Inst_3_U4  ( .A(\Red_MCInst_MC3_v1_2 [1]), .B(
        \MCInst_MC3_v1_0 [0]), .ZN(\MCInst_MC3_v1_2Inst_3_n3 ) );
  XOR2_X1 \MCInst_MC3_v1_2Inst_3_U3  ( .A(\MCInst_MC3_v1_3 [3]), .B(
        \Red_MCInst_MC3_v1_1 [2]), .Z(\MCInst_MC3_v1_2Inst_3_n4 ) );
  XOR2_X1 \MCInst_MC3_v2_1Inst_3_U3  ( .A(\MCInst_MC3_v2_0 [2]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\MCInst_MC3_v2_1 [3]) );
  XNOR2_X1 \MCInst_MC3_v2_2Inst_3_U4  ( .A(\MCInst_MC3_v2_2Inst_3_n2 ), .B(
        \MCInst_MC3_v2_0 [3]), .ZN(\MCInst_MC3_v2_2 [3]) );
  XNOR2_X1 \MCInst_MC3_v2_2Inst_3_U3  ( .A(\Red_MCInst_MC3_v2_2 [1]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\MCInst_MC3_v2_2Inst_3_n2 ) );
  XNOR2_X1 \MCInst_MC3_v2_3Inst_3_U4  ( .A(\MCInst_MC3_v2_3Inst_3_n2 ), .B(
        \MCInst_MC3_v2_0 [2]), .ZN(\MCInst_MC3_v2_3 [3]) );
  XNOR2_X1 \MCInst_MC3_v2_3Inst_3_U3  ( .A(\MCInst_MC3_v2_0 [3]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\MCInst_MC3_v2_3Inst_3_n2 ) );
  XOR2_X1 \MCInst_MC3_v3_1Inst_3_U3  ( .A(\Red_MCInst_MC3_v3_3 [2]), .B(
        \MCInst_MC3_v3_0 [3]), .Z(\MCInst_MC3_v3_1 [3]) );
  XOR2_X1 \MCInst_MC3_v3_3Inst_3_U3  ( .A(\MCInst_MC3_v3_2 [3]), .B(
        \MCInst_MC3_v3_0 [3]), .Z(\MCInst_MC3_v3_3 [3]) );
  XNOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC3_r0Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC3_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[48]) );
  XNOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_0_U2  ( .A(\Red_MCInst_MC3_v3_1 [2]), 
        .B(\Red_MCInst_MC3_v2_2 [1]), .ZN(\MCInst_MC3_r0Inst_XORInst_0_0_n4 )
         );
  XOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_0_U1  ( .A(\MCInst_MC3_v0_3 [3]), .B(
        \MCInst_MC3_v1_0 [0]), .Z(\MCInst_MC3_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC3_r0Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC3_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[49]) );
  XNOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_1_U2  ( .A(\MCInst_MC3_v3_0 [1]), .B(
        \MCInst_MC3_v2_0 [1]), .ZN(\MCInst_MC3_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_1_U1  ( .A(\MCInst_MC3_v0_0 [1]), .B(
        \Red_MCInst_MC3_v1_2 [1]), .Z(\MCInst_MC3_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC3_r0Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC3_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[50]) );
  XNOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_2_U2  ( .A(\Red_MCInst_MC3_v3_3 [2]), 
        .B(\MCInst_MC3_v2_0 [2]), .ZN(\MCInst_MC3_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_2_U1  ( .A(\MCInst_MC3_v0_0 [2]), .B(
        \MCInst_MC3_v1_3 [3]), .Z(\MCInst_MC3_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC3_r0Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC3_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[51]) );
  XNOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_3_U2  ( .A(\MCInst_MC3_v3_0 [3]), .B(
        \MCInst_MC3_v2_0 [3]), .ZN(\MCInst_MC3_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_3_U1  ( .A(\Red_MCInst_MC3_v0_2 [2]), 
        .B(\Red_MCInst_MC3_v1_1 [2]), .Z(\MCInst_MC3_r0Inst_XORInst_0_3_n5 )
         );
  XNOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC3_r1Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC3_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[32]) );
  XNOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_0_U2  ( .A(\MCInst_MC3_v3_1 [0]), .B(
        \MCInst_MC3_v2_1 [0]), .ZN(\MCInst_MC3_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC3_v0_2 [2]), 
        .B(\MCInst_MC3_v1_1 [0]), .Z(\MCInst_MC3_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC3_r1Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC3_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[33]) );
  XNOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_1_U2  ( .A(\MCInst_MC3_v3_1 [1]), .B(
        \MCInst_MC3_v2_1 [1]), .ZN(\MCInst_MC3_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_1_U1  ( .A(\MCInst_MC3_v0_1 [1]), .B(
        \MCInst_MC3_v1_1 [1]), .Z(\MCInst_MC3_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC3_r1Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC3_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[34]) );
  XNOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_2_U2  ( .A(\MCInst_MC3_v3_1 [2]), .B(
        \MCInst_MC3_v2_1 [2]), .ZN(\MCInst_MC3_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_2_U1  ( .A(\MCInst_MC3_v0_1 [2]), .B(
        \MCInst_MC3_v1_1 [2]), .Z(\MCInst_MC3_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC3_r1Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC3_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[35]) );
  XNOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_3_U2  ( .A(\MCInst_MC3_v3_1 [3]), .B(
        \MCInst_MC3_v2_1 [3]), .ZN(\MCInst_MC3_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_3_U1  ( .A(\MCInst_MC3_v0_1 [3]), .B(
        \MCInst_MC3_v1_1 [3]), .Z(\MCInst_MC3_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC3_r2Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC3_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[16]) );
  XNOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_0_U2  ( .A(\MCInst_MC3_v3_2 [0]), .B(
        \MCInst_MC3_v2_2 [0]), .ZN(\MCInst_MC3_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_0_U1  ( .A(\MCInst_MC3_v0_2 [0]), .B(
        \MCInst_MC3_v1_2 [0]), .Z(\MCInst_MC3_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC3_r2Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC3_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[17]) );
  XNOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_1_U2  ( .A(\MCInst_MC3_v3_0 [3]), .B(
        \MCInst_MC3_v2_2 [1]), .ZN(\MCInst_MC3_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_1_U1  ( .A(\MCInst_MC3_v0_2 [1]), .B(
        \MCInst_MC3_v1_2 [1]), .Z(\MCInst_MC3_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC3_r2Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC3_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[18]) );
  XNOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_2_U2  ( .A(\Red_MCInst_MC3_v3_1 [2]), 
        .B(\MCInst_MC3_v2_2 [2]), .ZN(\MCInst_MC3_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_2_U1  ( .A(\MCInst_MC3_v0_2 [2]), .B(
        \MCInst_MC3_v1_2 [2]), .Z(\MCInst_MC3_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC3_r2Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC3_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[19]) );
  XNOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_3_U2  ( .A(\MCInst_MC3_v3_2 [3]), .B(
        \MCInst_MC3_v2_2 [3]), .ZN(\MCInst_MC3_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_3_U1  ( .A(\MCInst_MC3_v0_2 [3]), .B(
        \MCInst_MC3_v1_2 [3]), .Z(\MCInst_MC3_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC3_r3Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC3_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[0]) );
  XNOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_0_U2  ( .A(\MCInst_MC3_v3_3 [0]), .B(
        \MCInst_MC3_v2_3 [0]), .ZN(\MCInst_MC3_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC3_v0_1 [0]), 
        .B(\Red_MCInst_MC3_v1_1 [2]), .Z(\MCInst_MC3_r3Inst_XORInst_0_0_n5 )
         );
  XNOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC3_r3Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC3_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[1]) );
  XNOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_1_U2  ( .A(\MCInst_MC3_v3_3 [1]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\MCInst_MC3_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_1_U1  ( .A(\MCInst_MC3_v0_3 [1]), .B(
        \MCInst_MC3_v1_3 [1]), .Z(\MCInst_MC3_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC3_r3Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC3_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[2]) );
  XNOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_2_U2  ( .A(\MCInst_MC3_v3_3 [2]), .B(
        \MCInst_MC3_v2_3 [2]), .ZN(\MCInst_MC3_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC3_v0_2 [2]), 
        .B(\Red_MCInst_MC3_v1_2 [1]), .Z(\MCInst_MC3_r3Inst_XORInst_0_2_n5 )
         );
  XNOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC3_r3Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC3_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[3]) );
  XNOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_3_U2  ( .A(\MCInst_MC3_v3_3 [3]), .B(
        \MCInst_MC3_v2_3 [3]), .ZN(\MCInst_MC3_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_3_U1  ( .A(\MCInst_MC3_v0_3 [3]), .B(
        \MCInst_MC3_v1_3 [3]), .Z(\MCInst_MC3_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_0_LFInst_0_n2 ), .B(Plaintext[1]), .ZN(
        Red_Plaintext[0]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_0_U3  ( .A(Plaintext[2]), .B(
        Plaintext[0]), .ZN(\Red_PlaintextInst_LFInst_0_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_0_LFInst_1_n2 ), .B(Plaintext[1]), .ZN(
        Red_Plaintext[1]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_1_U3  ( .A(Plaintext[3]), .B(
        Plaintext[0]), .ZN(\Red_PlaintextInst_LFInst_0_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_0_LFInst_2_n2 ), .B(Plaintext[2]), .ZN(
        Red_Plaintext[2]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_2_U3  ( .A(Plaintext[3]), .B(
        Plaintext[1]), .ZN(\Red_PlaintextInst_LFInst_0_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_1_LFInst_0_n2 ), .B(Plaintext[5]), .ZN(
        Red_Plaintext[3]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_0_U3  ( .A(Plaintext[6]), .B(
        Plaintext[4]), .ZN(\Red_PlaintextInst_LFInst_1_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_1_LFInst_1_n2 ), .B(Plaintext[5]), .ZN(
        Red_Plaintext[4]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_1_U3  ( .A(Plaintext[7]), .B(
        Plaintext[4]), .ZN(\Red_PlaintextInst_LFInst_1_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_1_LFInst_2_n2 ), .B(Plaintext[6]), .ZN(
        Red_Plaintext[5]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_2_U3  ( .A(Plaintext[7]), .B(
        Plaintext[5]), .ZN(\Red_PlaintextInst_LFInst_1_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_2_LFInst_0_n2 ), .B(Plaintext[9]), .ZN(
        Red_Plaintext[6]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_0_U3  ( .A(Plaintext[10]), .B(
        Plaintext[8]), .ZN(\Red_PlaintextInst_LFInst_2_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_2_LFInst_1_n2 ), .B(Plaintext[9]), .ZN(
        Red_Plaintext[7]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_1_U3  ( .A(Plaintext[11]), .B(
        Plaintext[8]), .ZN(\Red_PlaintextInst_LFInst_2_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_2_LFInst_2_n2 ), .B(Plaintext[10]), .ZN(
        Red_Plaintext[8]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_2_U3  ( .A(Plaintext[11]), .B(
        Plaintext[9]), .ZN(\Red_PlaintextInst_LFInst_2_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_3_LFInst_0_n2 ), .B(Plaintext[13]), .ZN(
        Red_Plaintext[9]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_0_U3  ( .A(Plaintext[14]), .B(
        Plaintext[12]), .ZN(\Red_PlaintextInst_LFInst_3_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_3_LFInst_1_n2 ), .B(Plaintext[13]), .ZN(
        Red_Plaintext[10]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_1_U3  ( .A(Plaintext[15]), .B(
        Plaintext[12]), .ZN(\Red_PlaintextInst_LFInst_3_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_3_LFInst_2_n2 ), .B(Plaintext[14]), .ZN(
        Red_Plaintext[11]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_2_U3  ( .A(Plaintext[15]), .B(
        Plaintext[13]), .ZN(\Red_PlaintextInst_LFInst_3_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_4_LFInst_0_n2 ), .B(Plaintext[17]), .ZN(
        Red_Plaintext[12]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_0_U3  ( .A(Plaintext[18]), .B(
        Plaintext[16]), .ZN(\Red_PlaintextInst_LFInst_4_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_4_LFInst_1_n2 ), .B(Plaintext[17]), .ZN(
        Red_Plaintext[13]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_1_U3  ( .A(Plaintext[19]), .B(
        Plaintext[16]), .ZN(\Red_PlaintextInst_LFInst_4_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_4_LFInst_2_n2 ), .B(Plaintext[18]), .ZN(
        Red_Plaintext[14]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_2_U3  ( .A(Plaintext[19]), .B(
        Plaintext[17]), .ZN(\Red_PlaintextInst_LFInst_4_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_5_LFInst_0_n2 ), .B(Plaintext[21]), .ZN(
        Red_Plaintext[15]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_0_U3  ( .A(Plaintext[22]), .B(
        Plaintext[20]), .ZN(\Red_PlaintextInst_LFInst_5_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_5_LFInst_1_n2 ), .B(Plaintext[21]), .ZN(
        Red_Plaintext[16]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_1_U3  ( .A(Plaintext[23]), .B(
        Plaintext[20]), .ZN(\Red_PlaintextInst_LFInst_5_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_5_LFInst_2_n2 ), .B(Plaintext[22]), .ZN(
        Red_Plaintext[17]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_2_U3  ( .A(Plaintext[23]), .B(
        Plaintext[21]), .ZN(\Red_PlaintextInst_LFInst_5_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_6_LFInst_0_n2 ), .B(Plaintext[25]), .ZN(
        Red_Plaintext[18]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_0_U3  ( .A(Plaintext[26]), .B(
        Plaintext[24]), .ZN(\Red_PlaintextInst_LFInst_6_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_6_LFInst_1_n2 ), .B(Plaintext[25]), .ZN(
        Red_Plaintext[19]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_1_U3  ( .A(Plaintext[27]), .B(
        Plaintext[24]), .ZN(\Red_PlaintextInst_LFInst_6_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_6_LFInst_2_n2 ), .B(Plaintext[26]), .ZN(
        Red_Plaintext[20]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_2_U3  ( .A(Plaintext[27]), .B(
        Plaintext[25]), .ZN(\Red_PlaintextInst_LFInst_6_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_7_LFInst_0_n2 ), .B(Plaintext[29]), .ZN(
        Red_Plaintext[21]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_0_U3  ( .A(Plaintext[30]), .B(
        Plaintext[28]), .ZN(\Red_PlaintextInst_LFInst_7_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_7_LFInst_1_n2 ), .B(Plaintext[29]), .ZN(
        Red_Plaintext[22]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_1_U3  ( .A(Plaintext[31]), .B(
        Plaintext[28]), .ZN(\Red_PlaintextInst_LFInst_7_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_7_LFInst_2_n2 ), .B(Plaintext[30]), .ZN(
        Red_Plaintext[23]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_2_U3  ( .A(Plaintext[31]), .B(
        Plaintext[29]), .ZN(\Red_PlaintextInst_LFInst_7_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_8_LFInst_0_n2 ), .B(Plaintext[33]), .ZN(
        Red_Plaintext[24]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_0_U3  ( .A(Plaintext[34]), .B(
        Plaintext[32]), .ZN(\Red_PlaintextInst_LFInst_8_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_8_LFInst_1_n2 ), .B(Plaintext[33]), .ZN(
        Red_Plaintext[25]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_1_U3  ( .A(Plaintext[35]), .B(
        Plaintext[32]), .ZN(\Red_PlaintextInst_LFInst_8_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_8_LFInst_2_n2 ), .B(Plaintext[34]), .ZN(
        Red_Plaintext[26]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_2_U3  ( .A(Plaintext[35]), .B(
        Plaintext[33]), .ZN(\Red_PlaintextInst_LFInst_8_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_9_LFInst_0_n2 ), .B(Plaintext[37]), .ZN(
        Red_Plaintext[27]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_0_U3  ( .A(Plaintext[38]), .B(
        Plaintext[36]), .ZN(\Red_PlaintextInst_LFInst_9_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_9_LFInst_1_n2 ), .B(Plaintext[37]), .ZN(
        Red_Plaintext[28]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_1_U3  ( .A(Plaintext[39]), .B(
        Plaintext[36]), .ZN(\Red_PlaintextInst_LFInst_9_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_9_LFInst_2_n2 ), .B(Plaintext[38]), .ZN(
        Red_Plaintext[29]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_2_U3  ( .A(Plaintext[39]), .B(
        Plaintext[37]), .ZN(\Red_PlaintextInst_LFInst_9_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_10_LFInst_0_n2 ), .B(Plaintext[41]), .ZN(
        Red_Plaintext[30]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_0_U3  ( .A(Plaintext[42]), .B(
        Plaintext[40]), .ZN(\Red_PlaintextInst_LFInst_10_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_10_LFInst_1_n2 ), .B(Plaintext[41]), .ZN(
        Red_Plaintext[31]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_1_U3  ( .A(Plaintext[43]), .B(
        Plaintext[40]), .ZN(\Red_PlaintextInst_LFInst_10_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_10_LFInst_2_n2 ), .B(Plaintext[42]), .ZN(
        Red_Plaintext[32]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_2_U3  ( .A(Plaintext[43]), .B(
        Plaintext[41]), .ZN(\Red_PlaintextInst_LFInst_10_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_11_LFInst_0_n2 ), .B(Plaintext[45]), .ZN(
        Red_Plaintext[33]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_0_U3  ( .A(Plaintext[46]), .B(
        Plaintext[44]), .ZN(\Red_PlaintextInst_LFInst_11_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_11_LFInst_1_n2 ), .B(Plaintext[45]), .ZN(
        Red_Plaintext[34]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_1_U3  ( .A(Plaintext[47]), .B(
        Plaintext[44]), .ZN(\Red_PlaintextInst_LFInst_11_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_11_LFInst_2_n2 ), .B(Plaintext[46]), .ZN(
        Red_Plaintext[35]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_2_U3  ( .A(Plaintext[47]), .B(
        Plaintext[45]), .ZN(\Red_PlaintextInst_LFInst_11_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_12_LFInst_0_n2 ), .B(Plaintext[49]), .ZN(
        Red_Plaintext[36]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_0_U3  ( .A(Plaintext[50]), .B(
        Plaintext[48]), .ZN(\Red_PlaintextInst_LFInst_12_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_12_LFInst_1_n2 ), .B(Plaintext[49]), .ZN(
        Red_Plaintext[37]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_1_U3  ( .A(Plaintext[51]), .B(
        Plaintext[48]), .ZN(\Red_PlaintextInst_LFInst_12_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_12_LFInst_2_n2 ), .B(Plaintext[50]), .ZN(
        Red_Plaintext[38]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_2_U3  ( .A(Plaintext[51]), .B(
        Plaintext[49]), .ZN(\Red_PlaintextInst_LFInst_12_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_13_LFInst_0_n2 ), .B(Plaintext[53]), .ZN(
        Red_Plaintext[39]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_0_U3  ( .A(Plaintext[54]), .B(
        Plaintext[52]), .ZN(\Red_PlaintextInst_LFInst_13_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_13_LFInst_1_n2 ), .B(Plaintext[53]), .ZN(
        Red_Plaintext[40]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_1_U3  ( .A(Plaintext[55]), .B(
        Plaintext[52]), .ZN(\Red_PlaintextInst_LFInst_13_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_13_LFInst_2_n2 ), .B(Plaintext[54]), .ZN(
        Red_Plaintext[41]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_2_U3  ( .A(Plaintext[55]), .B(
        Plaintext[53]), .ZN(\Red_PlaintextInst_LFInst_13_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_14_LFInst_0_n2 ), .B(Plaintext[57]), .ZN(
        Red_Plaintext[42]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_0_U3  ( .A(Plaintext[58]), .B(
        Plaintext[56]), .ZN(\Red_PlaintextInst_LFInst_14_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_14_LFInst_1_n2 ), .B(Plaintext[57]), .ZN(
        Red_Plaintext[43]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_1_U3  ( .A(Plaintext[59]), .B(
        Plaintext[56]), .ZN(\Red_PlaintextInst_LFInst_14_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_14_LFInst_2_n2 ), .B(Plaintext[58]), .ZN(
        Red_Plaintext[44]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_2_U3  ( .A(Plaintext[59]), .B(
        Plaintext[57]), .ZN(\Red_PlaintextInst_LFInst_14_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_15_LFInst_0_n2 ), .B(Plaintext[61]), .ZN(
        Red_Plaintext[45]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_0_U3  ( .A(Plaintext[62]), .B(
        Plaintext[60]), .ZN(\Red_PlaintextInst_LFInst_15_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_15_LFInst_1_n2 ), .B(Plaintext[61]), .ZN(
        Red_Plaintext[46]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_1_U3  ( .A(Plaintext[63]), .B(
        Plaintext[60]), .ZN(\Red_PlaintextInst_LFInst_15_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_15_LFInst_2_n2 ), .B(Plaintext[62]), .ZN(
        Red_Plaintext[47]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_2_U3  ( .A(Plaintext[63]), .B(
        Plaintext[61]), .ZN(\Red_PlaintextInst_LFInst_15_LFInst_2_n2 ) );
  DFF_X1 \Red_StateReg_s_current_state_reg[0]  ( .D(Red_Plaintext[0]), .CK(clk), .Q(Red_StateRegOutput[0]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[1]  ( .D(Red_Plaintext[1]), .CK(clk), .Q(Red_StateRegOutput[1]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[2]  ( .D(Red_Plaintext[2]), .CK(clk), .Q(Red_StateRegOutput[2]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[3]  ( .D(Red_Plaintext[3]), .CK(clk), .Q(Red_StateRegOutput[3]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[4]  ( .D(Red_Plaintext[4]), .CK(clk), .Q(Red_StateRegOutput[4]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[5]  ( .D(Red_Plaintext[5]), .CK(clk), .Q(Red_StateRegOutput[5]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[6]  ( .D(Red_Plaintext[6]), .CK(clk), .Q(Red_AddConstOutput[0]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[7]  ( .D(Red_Plaintext[7]), .CK(clk), .Q(Red_AddConstOutput[1]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[8]  ( .D(Red_Plaintext[8]), .CK(clk), .Q(Red_AddConstOutput[2]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[9]  ( .D(Red_Plaintext[9]), .CK(clk), .Q(Red_AddConstOutput[3]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[10]  ( .D(Red_Plaintext[10]), .CK(
        clk), .Q(Red_AddConstOutput[4]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[11]  ( .D(Red_Plaintext[11]), .CK(
        clk), .Q(Red_StateRegOutput[11]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[12]  ( .D(Red_Plaintext[12]), .CK(
        clk), .Q(Red_StateRegOutput[12]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[13]  ( .D(Red_Plaintext[13]), .CK(
        clk), .Q(Red_StateRegOutput[13]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[14]  ( .D(Red_Plaintext[14]), .CK(
        clk), .Q(Red_StateRegOutput[14]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[15]  ( .D(Red_Plaintext[15]), .CK(
        clk), .Q(Red_StateRegOutput[15]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[16]  ( .D(Red_Plaintext[16]), .CK(
        clk), .Q(Red_StateRegOutput[16]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[17]  ( .D(Red_Plaintext[17]), .CK(
        clk), .Q(Red_StateRegOutput[17]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[18]  ( .D(Red_Plaintext[18]), .CK(
        clk), .Q(Red_AddConstOutput[6]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[19]  ( .D(Red_Plaintext[19]), .CK(
        clk), .Q(Red_AddConstOutput[7]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[20]  ( .D(Red_Plaintext[20]), .CK(
        clk), .Q(Red_AddConstOutput[8]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[21]  ( .D(Red_Plaintext[21]), .CK(
        clk), .Q(Red_StateRegOutput[21]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[22]  ( .D(Red_Plaintext[22]), .CK(
        clk), .Q(Red_StateRegOutput[22]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[23]  ( .D(Red_Plaintext[23]), .CK(
        clk), .Q(Red_StateRegOutput[23]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[24]  ( .D(Red_Plaintext[24]), .CK(
        clk), .Q(Red_StateRegOutput[24]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[25]  ( .D(Red_Plaintext[25]), .CK(
        clk), .Q(Red_StateRegOutput[25]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[26]  ( .D(Red_Plaintext[26]), .CK(
        clk), .Q(Red_StateRegOutput[26]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[27]  ( .D(Red_Plaintext[27]), .CK(
        clk), .Q(Red_StateRegOutput[27]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[28]  ( .D(Red_Plaintext[28]), .CK(
        clk), .Q(Red_StateRegOutput[28]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[29]  ( .D(Red_Plaintext[29]), .CK(
        clk), .Q(Red_StateRegOutput[29]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[30]  ( .D(Red_Plaintext[30]), .CK(
        clk), .Q(Red_AddConstOutput[12]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[31]  ( .D(Red_Plaintext[31]), .CK(
        clk), .Q(Red_AddConstOutput[13]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[32]  ( .D(Red_Plaintext[32]), .CK(
        clk), .Q(Red_AddConstOutput[14]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[33]  ( .D(Red_Plaintext[33]), .CK(
        clk), .Q(Red_AddConstOutput[15]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[34]  ( .D(Red_Plaintext[34]), .CK(
        clk), .Q(Red_StateRegOutput[34]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[35]  ( .D(Red_Plaintext[35]), .CK(
        clk), .Q(Red_StateRegOutput[35]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[36]  ( .D(Red_Plaintext[36]), .CK(
        clk), .Q(Red_StateRegOutput[36]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[37]  ( .D(Red_Plaintext[37]), .CK(
        clk), .Q(Red_StateRegOutput[37]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[38]  ( .D(Red_Plaintext[38]), .CK(
        clk), .Q(Red_StateRegOutput[38]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[39]  ( .D(Red_Plaintext[39]), .CK(
        clk), .Q(Red_StateRegOutput[39]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[40]  ( .D(Red_Plaintext[40]), .CK(
        clk), .Q(Red_StateRegOutput[40]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[41]  ( .D(Red_Plaintext[41]), .CK(
        clk), .Q(Red_StateRegOutput[41]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[42]  ( .D(Red_Plaintext[42]), .CK(
        clk), .Q(Red_AddConstOutput[18]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[43]  ( .D(Red_Plaintext[43]), .CK(
        clk), .Q(Red_AddConstOutput[19]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[44]  ( .D(Red_Plaintext[44]), .CK(
        clk), .Q(Red_AddConstOutput[20]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[45]  ( .D(Red_Plaintext[45]), .CK(
        clk), .Q(Red_StateRegOutput[45]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[46]  ( .D(Red_Plaintext[46]), .CK(
        clk), .Q(Red_AddConstOutput[22]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[47]  ( .D(Red_Plaintext[47]), .CK(
        clk), .Q(Red_StateRegOutput[47]) );
  INV_X1 \Red_AddConstXOR_XORInst_XORInst_1_2_U1  ( .A(Red_StateRegOutput[11]), 
        .ZN(Red_AddConstOutput[5]) );
  INV_X1 \Red_AddConstXOR_XORInst_XORInst_3_0_U1  ( .A(Red_StateRegOutput[21]), 
        .ZN(Red_AddConstOutput[9]) );
  INV_X1 \Red_AddConstXOR_XORInst_XORInst_3_1_U1  ( .A(Red_StateRegOutput[22]), 
        .ZN(Red_AddConstOutput[10]) );
  INV_X1 \Red_AddConstXOR_XORInst_XORInst_3_2_U1  ( .A(Red_StateRegOutput[23]), 
        .ZN(Red_AddConstOutput[11]) );
  INV_X1 \Red_AddConstXOR_XORInst_XORInst_5_1_U1  ( .A(Red_StateRegOutput[34]), 
        .ZN(Red_AddConstOutput[16]) );
  INV_X1 \Red_AddConstXOR_XORInst_XORInst_5_2_U1  ( .A(Red_StateRegOutput[35]), 
        .ZN(Red_AddConstOutput[17]) );
  INV_X1 \Red_AddConstXOR_XORInst_XORInst_7_0_U1  ( .A(Red_StateRegOutput[45]), 
        .ZN(Red_AddConstOutput[21]) );
  INV_X1 \Red_AddConstXOR_XORInst_XORInst_7_2_U1  ( .A(Red_StateRegOutput[47]), 
        .ZN(Red_AddConstOutput[23]) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U7  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_0_n8 ), .A2(
        \Red_SubCellInst_LFInst_0_LFInst_0_n7 ), .ZN(Red_ShiftRowsOutput[9])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U6  ( .A1(StateRegOutput[2]), 
        .A2(StateRegOutput[3]), .ZN(\Red_SubCellInst_LFInst_0_LFInst_0_n7 ) );
  OR2_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U5  ( .A1(StateRegOutput[0]), .A2(
        \Red_SubCellInst_LFInst_0_LFInst_0_n6 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_0_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U4  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_0_n5 ), .A2(StateRegOutput[2]), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_0_n6 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U3  ( .A(StateRegOutput[1]), .B(
        StateRegOutput[3]), .ZN(\Red_SubCellInst_LFInst_0_LFInst_0_n5 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_1_U5  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_1_n4 ), .A2(
        \Red_SubCellInst_LFInst_0_LFInst_1_n3 ), .ZN(Red_ShiftRowsOutput[10])
         );
  OR2_X1 \Red_SubCellInst_LFInst_0_LFInst_1_U4  ( .A1(StateRegOutput[3]), .A2(
        StateRegOutput[2]), .ZN(\Red_SubCellInst_LFInst_0_LFInst_1_n3 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_1_U3  ( .A1(StateRegOutput[1]), 
        .A2(StateRegOutput[3]), .ZN(\Red_SubCellInst_LFInst_0_LFInst_1_n4 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U8  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_2_n11 ), .A2(
        \Red_SubCellInst_LFInst_0_LFInst_2_n10 ), .ZN(Red_ShiftRowsOutput[11])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U7  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_2_n9 ), .A2(StateRegOutput[3]), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_2_n10 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U6  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_2_n8 ), .A2(StateRegOutput[2]), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_2_n9 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U5  ( .A1(StateRegOutput[0]), 
        .A2(StateRegOutput[1]), .ZN(\Red_SubCellInst_LFInst_0_LFInst_2_n8 ) );
  OR2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U4  ( .A1(StateRegOutput[1]), .A2(
        \Red_SubCellInst_LFInst_0_LFInst_2_n7 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_2_n11 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U3  ( .A(StateRegOutput[2]), .B(
        StateRegOutput[0]), .ZN(\Red_SubCellInst_LFInst_0_LFInst_2_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U7  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_0_n8 ), .A2(
        \Red_SubCellInst_LFInst_1_LFInst_0_n7 ), .ZN(Red_ShiftRowsOutput[0])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U6  ( .A1(StateRegOutput[6]), 
        .A2(StateRegOutput[7]), .ZN(\Red_SubCellInst_LFInst_1_LFInst_0_n7 ) );
  OR2_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U5  ( .A1(StateRegOutput[4]), .A2(
        \Red_SubCellInst_LFInst_1_LFInst_0_n6 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_0_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U4  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_0_n5 ), .A2(StateRegOutput[6]), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_0_n6 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U3  ( .A(StateRegOutput[5]), .B(
        StateRegOutput[7]), .ZN(\Red_SubCellInst_LFInst_1_LFInst_0_n5 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_1_U5  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_1_n4 ), .A2(
        \Red_SubCellInst_LFInst_1_LFInst_1_n3 ), .ZN(Red_ShiftRowsOutput[1])
         );
  OR2_X1 \Red_SubCellInst_LFInst_1_LFInst_1_U4  ( .A1(StateRegOutput[7]), .A2(
        StateRegOutput[6]), .ZN(\Red_SubCellInst_LFInst_1_LFInst_1_n3 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_1_U3  ( .A1(StateRegOutput[5]), 
        .A2(StateRegOutput[7]), .ZN(\Red_SubCellInst_LFInst_1_LFInst_1_n4 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U8  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_2_n11 ), .A2(
        \Red_SubCellInst_LFInst_1_LFInst_2_n10 ), .ZN(Red_ShiftRowsOutput[2])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U7  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_2_n9 ), .A2(StateRegOutput[7]), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_2_n10 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U6  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_2_n8 ), .A2(StateRegOutput[6]), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_2_n9 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U5  ( .A1(StateRegOutput[4]), 
        .A2(StateRegOutput[5]), .ZN(\Red_SubCellInst_LFInst_1_LFInst_2_n8 ) );
  OR2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U4  ( .A1(StateRegOutput[5]), .A2(
        \Red_SubCellInst_LFInst_1_LFInst_2_n7 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_2_n11 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U3  ( .A(StateRegOutput[6]), .B(
        StateRegOutput[4]), .ZN(\Red_SubCellInst_LFInst_1_LFInst_2_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U7  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_0_n8 ), .A2(
        \Red_SubCellInst_LFInst_2_LFInst_0_n7 ), .ZN(Red_ShiftRowsOutput[3])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U6  ( .A1(AddConstOutput[2]), 
        .A2(AddConstOutput[3]), .ZN(\Red_SubCellInst_LFInst_2_LFInst_0_n7 ) );
  OR2_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U5  ( .A1(AddConstOutput[0]), .A2(
        \Red_SubCellInst_LFInst_2_LFInst_0_n6 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_0_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U4  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_0_n5 ), .A2(AddConstOutput[2]), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_0_n6 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U3  ( .A(AddConstOutput[1]), .B(
        AddConstOutput[3]), .ZN(\Red_SubCellInst_LFInst_2_LFInst_0_n5 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_1_U5  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_1_n4 ), .A2(
        \Red_SubCellInst_LFInst_2_LFInst_1_n3 ), .ZN(Red_ShiftRowsOutput[4])
         );
  OR2_X1 \Red_SubCellInst_LFInst_2_LFInst_1_U4  ( .A1(AddConstOutput[3]), .A2(
        AddConstOutput[2]), .ZN(\Red_SubCellInst_LFInst_2_LFInst_1_n3 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_1_U3  ( .A1(AddConstOutput[1]), 
        .A2(AddConstOutput[3]), .ZN(\Red_SubCellInst_LFInst_2_LFInst_1_n4 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U8  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_2_n11 ), .A2(
        \Red_SubCellInst_LFInst_2_LFInst_2_n10 ), .ZN(Red_ShiftRowsOutput[5])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U7  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_2_n9 ), .A2(AddConstOutput[3]), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_2_n10 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U6  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_2_n8 ), .A2(AddConstOutput[2]), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_2_n9 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U5  ( .A1(AddConstOutput[0]), 
        .A2(AddConstOutput[1]), .ZN(\Red_SubCellInst_LFInst_2_LFInst_2_n8 ) );
  OR2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U4  ( .A1(AddConstOutput[1]), .A2(
        \Red_SubCellInst_LFInst_2_LFInst_2_n7 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_2_n11 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U3  ( .A(AddConstOutput[2]), .B(
        AddConstOutput[0]), .ZN(\Red_SubCellInst_LFInst_2_LFInst_2_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U7  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_0_n8 ), .A2(
        \Red_SubCellInst_LFInst_3_LFInst_0_n7 ), .ZN(Red_ShiftRowsOutput[6])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U6  ( .A1(AddConstOutput[6]), 
        .A2(AddConstOutput[7]), .ZN(\Red_SubCellInst_LFInst_3_LFInst_0_n7 ) );
  OR2_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U5  ( .A1(AddConstOutput[4]), .A2(
        \Red_SubCellInst_LFInst_3_LFInst_0_n6 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_0_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U4  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_0_n5 ), .A2(AddConstOutput[6]), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_0_n6 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U3  ( .A(AddConstOutput[5]), .B(
        AddConstOutput[7]), .ZN(\Red_SubCellInst_LFInst_3_LFInst_0_n5 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_1_U5  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_1_n4 ), .A2(
        \Red_SubCellInst_LFInst_3_LFInst_1_n3 ), .ZN(Red_ShiftRowsOutput[7])
         );
  OR2_X1 \Red_SubCellInst_LFInst_3_LFInst_1_U4  ( .A1(AddConstOutput[7]), .A2(
        AddConstOutput[6]), .ZN(\Red_SubCellInst_LFInst_3_LFInst_1_n3 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_1_U3  ( .A1(AddConstOutput[5]), 
        .A2(AddConstOutput[7]), .ZN(\Red_SubCellInst_LFInst_3_LFInst_1_n4 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U8  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_2_n11 ), .A2(
        \Red_SubCellInst_LFInst_3_LFInst_2_n10 ), .ZN(Red_ShiftRowsOutput[8])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U7  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_2_n9 ), .A2(AddConstOutput[7]), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_2_n10 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U6  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_2_n8 ), .A2(AddConstOutput[6]), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_2_n9 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U5  ( .A1(AddConstOutput[4]), 
        .A2(AddConstOutput[5]), .ZN(\Red_SubCellInst_LFInst_3_LFInst_2_n8 ) );
  OR2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U4  ( .A1(AddConstOutput[5]), .A2(
        \Red_SubCellInst_LFInst_3_LFInst_2_n7 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_2_n11 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U3  ( .A(AddConstOutput[6]), .B(
        AddConstOutput[4]), .ZN(\Red_SubCellInst_LFInst_3_LFInst_2_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U7  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_0_n8 ), .A2(
        \Red_SubCellInst_LFInst_4_LFInst_0_n7 ), .ZN(Red_ShiftRowsOutput[18])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U6  ( .A1(StateRegOutput[18]), 
        .A2(StateRegOutput[19]), .ZN(\Red_SubCellInst_LFInst_4_LFInst_0_n7 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U5  ( .A1(StateRegOutput[16]), 
        .A2(\Red_SubCellInst_LFInst_4_LFInst_0_n6 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_0_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U4  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_0_n5 ), .A2(StateRegOutput[18]), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_0_n6 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U3  ( .A(StateRegOutput[17]), 
        .B(StateRegOutput[19]), .ZN(\Red_SubCellInst_LFInst_4_LFInst_0_n5 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_1_U5  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_1_n4 ), .A2(
        \Red_SubCellInst_LFInst_4_LFInst_1_n3 ), .ZN(Red_ShiftRowsOutput[19])
         );
  OR2_X1 \Red_SubCellInst_LFInst_4_LFInst_1_U4  ( .A1(StateRegOutput[19]), 
        .A2(StateRegOutput[18]), .ZN(\Red_SubCellInst_LFInst_4_LFInst_1_n3 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_1_U3  ( .A1(StateRegOutput[17]), 
        .A2(StateRegOutput[19]), .ZN(\Red_SubCellInst_LFInst_4_LFInst_1_n4 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U8  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_2_n11 ), .A2(
        \Red_SubCellInst_LFInst_4_LFInst_2_n10 ), .ZN(Red_ShiftRowsOutput[20])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U7  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_2_n9 ), .A2(StateRegOutput[19]), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_2_n10 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U6  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_2_n8 ), .A2(StateRegOutput[18]), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_2_n9 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U5  ( .A1(StateRegOutput[16]), 
        .A2(StateRegOutput[17]), .ZN(\Red_SubCellInst_LFInst_4_LFInst_2_n8 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U4  ( .A1(StateRegOutput[17]), 
        .A2(\Red_SubCellInst_LFInst_4_LFInst_2_n7 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_2_n11 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U3  ( .A(StateRegOutput[18]), 
        .B(StateRegOutput[16]), .ZN(\Red_SubCellInst_LFInst_4_LFInst_2_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U7  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_0_n8 ), .A2(
        \Red_SubCellInst_LFInst_5_LFInst_0_n7 ), .ZN(Red_ShiftRowsOutput[21])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U6  ( .A1(StateRegOutput[22]), 
        .A2(StateRegOutput[23]), .ZN(\Red_SubCellInst_LFInst_5_LFInst_0_n7 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U5  ( .A1(StateRegOutput[20]), 
        .A2(\Red_SubCellInst_LFInst_5_LFInst_0_n6 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_0_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U4  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_0_n5 ), .A2(StateRegOutput[22]), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_0_n6 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U3  ( .A(StateRegOutput[21]), 
        .B(StateRegOutput[23]), .ZN(\Red_SubCellInst_LFInst_5_LFInst_0_n5 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_1_U5  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_1_n4 ), .A2(
        \Red_SubCellInst_LFInst_5_LFInst_1_n3 ), .ZN(Red_ShiftRowsOutput[22])
         );
  OR2_X1 \Red_SubCellInst_LFInst_5_LFInst_1_U4  ( .A1(StateRegOutput[23]), 
        .A2(StateRegOutput[22]), .ZN(\Red_SubCellInst_LFInst_5_LFInst_1_n3 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_1_U3  ( .A1(StateRegOutput[21]), 
        .A2(StateRegOutput[23]), .ZN(\Red_SubCellInst_LFInst_5_LFInst_1_n4 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U8  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_2_n11 ), .A2(
        \Red_SubCellInst_LFInst_5_LFInst_2_n10 ), .ZN(Red_ShiftRowsOutput[23])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U7  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_2_n9 ), .A2(StateRegOutput[23]), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_2_n10 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U6  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_2_n8 ), .A2(StateRegOutput[22]), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_2_n9 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U5  ( .A1(StateRegOutput[20]), 
        .A2(StateRegOutput[21]), .ZN(\Red_SubCellInst_LFInst_5_LFInst_2_n8 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U4  ( .A1(StateRegOutput[21]), 
        .A2(\Red_SubCellInst_LFInst_5_LFInst_2_n7 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_2_n11 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U3  ( .A(StateRegOutput[22]), 
        .B(StateRegOutput[20]), .ZN(\Red_SubCellInst_LFInst_5_LFInst_2_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U7  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_0_n8 ), .A2(
        \Red_SubCellInst_LFInst_6_LFInst_0_n7 ), .ZN(Red_ShiftRowsOutput[12])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U6  ( .A1(AddConstOutput[10]), 
        .A2(AddConstOutput[11]), .ZN(\Red_SubCellInst_LFInst_6_LFInst_0_n7 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U5  ( .A1(AddConstOutput[8]), .A2(
        \Red_SubCellInst_LFInst_6_LFInst_0_n6 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_0_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U4  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_0_n5 ), .A2(AddConstOutput[10]), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_0_n6 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U3  ( .A(AddConstOutput[9]), .B(
        AddConstOutput[11]), .ZN(\Red_SubCellInst_LFInst_6_LFInst_0_n5 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_1_U5  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_1_n4 ), .A2(
        \Red_SubCellInst_LFInst_6_LFInst_1_n3 ), .ZN(Red_ShiftRowsOutput[13])
         );
  OR2_X1 \Red_SubCellInst_LFInst_6_LFInst_1_U4  ( .A1(AddConstOutput[11]), 
        .A2(AddConstOutput[10]), .ZN(\Red_SubCellInst_LFInst_6_LFInst_1_n3 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_1_U3  ( .A1(AddConstOutput[9]), 
        .A2(AddConstOutput[11]), .ZN(\Red_SubCellInst_LFInst_6_LFInst_1_n4 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U8  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_2_n11 ), .A2(
        \Red_SubCellInst_LFInst_6_LFInst_2_n10 ), .ZN(Red_ShiftRowsOutput[14])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U7  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_2_n9 ), .A2(AddConstOutput[11]), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_2_n10 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U6  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_2_n8 ), .A2(AddConstOutput[10]), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_2_n9 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U5  ( .A1(AddConstOutput[8]), 
        .A2(AddConstOutput[9]), .ZN(\Red_SubCellInst_LFInst_6_LFInst_2_n8 ) );
  OR2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U4  ( .A1(AddConstOutput[9]), .A2(
        \Red_SubCellInst_LFInst_6_LFInst_2_n7 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_2_n11 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U3  ( .A(AddConstOutput[10]), 
        .B(AddConstOutput[8]), .ZN(\Red_SubCellInst_LFInst_6_LFInst_2_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U7  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_0_n8 ), .A2(
        \Red_SubCellInst_LFInst_7_LFInst_0_n7 ), .ZN(Red_ShiftRowsOutput[15])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U6  ( .A1(AddConstOutput[14]), 
        .A2(AddConstOutput[15]), .ZN(\Red_SubCellInst_LFInst_7_LFInst_0_n7 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U5  ( .A1(AddConstOutput[12]), 
        .A2(\Red_SubCellInst_LFInst_7_LFInst_0_n6 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_0_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U4  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_0_n5 ), .A2(AddConstOutput[14]), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_0_n6 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U3  ( .A(AddConstOutput[13]), 
        .B(AddConstOutput[15]), .ZN(\Red_SubCellInst_LFInst_7_LFInst_0_n5 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_1_U5  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_1_n4 ), .A2(
        \Red_SubCellInst_LFInst_7_LFInst_1_n3 ), .ZN(Red_ShiftRowsOutput[16])
         );
  OR2_X1 \Red_SubCellInst_LFInst_7_LFInst_1_U4  ( .A1(AddConstOutput[15]), 
        .A2(AddConstOutput[14]), .ZN(\Red_SubCellInst_LFInst_7_LFInst_1_n3 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_1_U3  ( .A1(AddConstOutput[13]), 
        .A2(AddConstOutput[15]), .ZN(\Red_SubCellInst_LFInst_7_LFInst_1_n4 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U8  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_2_n11 ), .A2(
        \Red_SubCellInst_LFInst_7_LFInst_2_n10 ), .ZN(Red_ShiftRowsOutput[17])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U7  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_2_n9 ), .A2(AddConstOutput[15]), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_2_n10 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U6  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_2_n8 ), .A2(AddConstOutput[14]), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_2_n9 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U5  ( .A1(AddConstOutput[12]), 
        .A2(AddConstOutput[13]), .ZN(\Red_SubCellInst_LFInst_7_LFInst_2_n8 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U4  ( .A1(AddConstOutput[13]), 
        .A2(\Red_SubCellInst_LFInst_7_LFInst_2_n7 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_2_n11 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U3  ( .A(AddConstOutput[14]), 
        .B(AddConstOutput[12]), .ZN(\Red_SubCellInst_LFInst_7_LFInst_2_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U7  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_0_n8 ), .A2(
        \Red_SubCellInst_LFInst_8_LFInst_0_n7 ), .ZN(Red_ShiftRowsOutput[27])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U6  ( .A1(StateRegOutput[34]), 
        .A2(StateRegOutput[35]), .ZN(\Red_SubCellInst_LFInst_8_LFInst_0_n7 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U5  ( .A1(StateRegOutput[32]), 
        .A2(\Red_SubCellInst_LFInst_8_LFInst_0_n6 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_0_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U4  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_0_n5 ), .A2(StateRegOutput[34]), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_0_n6 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U3  ( .A(StateRegOutput[33]), 
        .B(StateRegOutput[35]), .ZN(\Red_SubCellInst_LFInst_8_LFInst_0_n5 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_1_U5  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_1_n4 ), .A2(
        \Red_SubCellInst_LFInst_8_LFInst_1_n3 ), .ZN(Red_ShiftRowsOutput[28])
         );
  OR2_X1 \Red_SubCellInst_LFInst_8_LFInst_1_U4  ( .A1(StateRegOutput[35]), 
        .A2(StateRegOutput[34]), .ZN(\Red_SubCellInst_LFInst_8_LFInst_1_n3 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_1_U3  ( .A1(StateRegOutput[33]), 
        .A2(StateRegOutput[35]), .ZN(\Red_SubCellInst_LFInst_8_LFInst_1_n4 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U8  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_2_n11 ), .A2(
        \Red_SubCellInst_LFInst_8_LFInst_2_n10 ), .ZN(Red_ShiftRowsOutput[29])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U7  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_2_n9 ), .A2(StateRegOutput[35]), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_2_n10 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U6  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_2_n8 ), .A2(StateRegOutput[34]), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_2_n9 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U5  ( .A1(StateRegOutput[32]), 
        .A2(StateRegOutput[33]), .ZN(\Red_SubCellInst_LFInst_8_LFInst_2_n8 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U4  ( .A1(StateRegOutput[33]), 
        .A2(\Red_SubCellInst_LFInst_8_LFInst_2_n7 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_2_n11 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U3  ( .A(StateRegOutput[34]), 
        .B(StateRegOutput[32]), .ZN(\Red_SubCellInst_LFInst_8_LFInst_2_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U7  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_0_n8 ), .A2(
        \Red_SubCellInst_LFInst_9_LFInst_0_n7 ), .ZN(Red_ShiftRowsOutput[30])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U6  ( .A1(StateRegOutput[38]), 
        .A2(StateRegOutput[39]), .ZN(\Red_SubCellInst_LFInst_9_LFInst_0_n7 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U5  ( .A1(StateRegOutput[36]), 
        .A2(\Red_SubCellInst_LFInst_9_LFInst_0_n6 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_0_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U4  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_0_n5 ), .A2(StateRegOutput[38]), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_0_n6 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U3  ( .A(StateRegOutput[37]), 
        .B(StateRegOutput[39]), .ZN(\Red_SubCellInst_LFInst_9_LFInst_0_n5 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_1_U5  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_1_n4 ), .A2(
        \Red_SubCellInst_LFInst_9_LFInst_1_n3 ), .ZN(Red_ShiftRowsOutput[31])
         );
  OR2_X1 \Red_SubCellInst_LFInst_9_LFInst_1_U4  ( .A1(StateRegOutput[39]), 
        .A2(StateRegOutput[38]), .ZN(\Red_SubCellInst_LFInst_9_LFInst_1_n3 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_1_U3  ( .A1(StateRegOutput[37]), 
        .A2(StateRegOutput[39]), .ZN(\Red_SubCellInst_LFInst_9_LFInst_1_n4 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U8  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_2_n11 ), .A2(
        \Red_SubCellInst_LFInst_9_LFInst_2_n10 ), .ZN(Red_ShiftRowsOutput[32])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U7  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_2_n9 ), .A2(StateRegOutput[39]), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_2_n10 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U6  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_2_n8 ), .A2(StateRegOutput[38]), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_2_n9 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U5  ( .A1(StateRegOutput[36]), 
        .A2(StateRegOutput[37]), .ZN(\Red_SubCellInst_LFInst_9_LFInst_2_n8 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U4  ( .A1(StateRegOutput[37]), 
        .A2(\Red_SubCellInst_LFInst_9_LFInst_2_n7 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_2_n11 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U3  ( .A(StateRegOutput[38]), 
        .B(StateRegOutput[36]), .ZN(\Red_SubCellInst_LFInst_9_LFInst_2_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U7  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_0_n8 ), .A2(
        \Red_SubCellInst_LFInst_10_LFInst_0_n7 ), .ZN(Red_ShiftRowsOutput[33])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U6  ( .A1(AddConstOutput[18]), 
        .A2(AddConstOutput[19]), .ZN(\Red_SubCellInst_LFInst_10_LFInst_0_n7 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U5  ( .A1(AddConstOutput[16]), 
        .A2(\Red_SubCellInst_LFInst_10_LFInst_0_n6 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_0_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U4  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_0_n5 ), .A2(AddConstOutput[18]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_0_n6 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U3  ( .A(AddConstOutput[17]), 
        .B(AddConstOutput[19]), .ZN(\Red_SubCellInst_LFInst_10_LFInst_0_n5 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_1_U5  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_1_n4 ), .A2(
        \Red_SubCellInst_LFInst_10_LFInst_1_n3 ), .ZN(Red_ShiftRowsOutput[34])
         );
  OR2_X1 \Red_SubCellInst_LFInst_10_LFInst_1_U4  ( .A1(AddConstOutput[19]), 
        .A2(AddConstOutput[18]), .ZN(\Red_SubCellInst_LFInst_10_LFInst_1_n3 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_1_U3  ( .A1(AddConstOutput[17]), 
        .A2(AddConstOutput[19]), .ZN(\Red_SubCellInst_LFInst_10_LFInst_1_n4 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U8  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_2_n11 ), .A2(
        \Red_SubCellInst_LFInst_10_LFInst_2_n10 ), .ZN(Red_ShiftRowsOutput[35]) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U7  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_2_n9 ), .A2(AddConstOutput[19]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_2_n10 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U6  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_2_n8 ), .A2(AddConstOutput[18]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_2_n9 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U5  ( .A1(AddConstOutput[16]), 
        .A2(AddConstOutput[17]), .ZN(\Red_SubCellInst_LFInst_10_LFInst_2_n8 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U4  ( .A1(AddConstOutput[17]), 
        .A2(\Red_SubCellInst_LFInst_10_LFInst_2_n7 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_2_n11 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U3  ( .A(AddConstOutput[18]), 
        .B(AddConstOutput[16]), .ZN(\Red_SubCellInst_LFInst_10_LFInst_2_n7 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U7  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_0_n8 ), .A2(
        \Red_SubCellInst_LFInst_11_LFInst_0_n7 ), .ZN(Red_ShiftRowsOutput[24])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U6  ( .A1(AddConstOutput[22]), 
        .A2(AddConstOutput[23]), .ZN(\Red_SubCellInst_LFInst_11_LFInst_0_n7 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U5  ( .A1(AddConstOutput[20]), 
        .A2(\Red_SubCellInst_LFInst_11_LFInst_0_n6 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_0_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U4  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_0_n5 ), .A2(AddConstOutput[22]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_0_n6 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U3  ( .A(AddConstOutput[21]), 
        .B(AddConstOutput[23]), .ZN(\Red_SubCellInst_LFInst_11_LFInst_0_n5 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_1_U5  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_1_n4 ), .A2(
        \Red_SubCellInst_LFInst_11_LFInst_1_n3 ), .ZN(Red_ShiftRowsOutput[25])
         );
  OR2_X1 \Red_SubCellInst_LFInst_11_LFInst_1_U4  ( .A1(AddConstOutput[23]), 
        .A2(AddConstOutput[22]), .ZN(\Red_SubCellInst_LFInst_11_LFInst_1_n3 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_1_U3  ( .A1(AddConstOutput[21]), 
        .A2(AddConstOutput[23]), .ZN(\Red_SubCellInst_LFInst_11_LFInst_1_n4 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U8  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_2_n11 ), .A2(
        \Red_SubCellInst_LFInst_11_LFInst_2_n10 ), .ZN(Red_ShiftRowsOutput[26]) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U7  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_2_n9 ), .A2(AddConstOutput[23]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_2_n10 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U6  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_2_n8 ), .A2(AddConstOutput[22]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_2_n9 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U5  ( .A1(AddConstOutput[20]), 
        .A2(AddConstOutput[21]), .ZN(\Red_SubCellInst_LFInst_11_LFInst_2_n8 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U4  ( .A1(AddConstOutput[21]), 
        .A2(\Red_SubCellInst_LFInst_11_LFInst_2_n7 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_2_n11 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U3  ( .A(AddConstOutput[22]), 
        .B(AddConstOutput[20]), .ZN(\Red_SubCellInst_LFInst_11_LFInst_2_n7 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U7  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_0_n8 ), .A2(
        \Red_SubCellInst_LFInst_12_LFInst_0_n7 ), .ZN(Red_ShiftRowsOutput[36])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U6  ( .A1(StateRegOutput[50]), 
        .A2(StateRegOutput[51]), .ZN(\Red_SubCellInst_LFInst_12_LFInst_0_n7 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U5  ( .A1(StateRegOutput[48]), 
        .A2(\Red_SubCellInst_LFInst_12_LFInst_0_n6 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_0_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U4  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_0_n5 ), .A2(StateRegOutput[50]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_0_n6 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U3  ( .A(StateRegOutput[49]), 
        .B(StateRegOutput[51]), .ZN(\Red_SubCellInst_LFInst_12_LFInst_0_n5 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_1_U5  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_1_n4 ), .A2(
        \Red_SubCellInst_LFInst_12_LFInst_1_n3 ), .ZN(Red_ShiftRowsOutput[37])
         );
  OR2_X1 \Red_SubCellInst_LFInst_12_LFInst_1_U4  ( .A1(StateRegOutput[51]), 
        .A2(StateRegOutput[50]), .ZN(\Red_SubCellInst_LFInst_12_LFInst_1_n3 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_1_U3  ( .A1(StateRegOutput[49]), 
        .A2(StateRegOutput[51]), .ZN(\Red_SubCellInst_LFInst_12_LFInst_1_n4 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U8  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_2_n11 ), .A2(
        \Red_SubCellInst_LFInst_12_LFInst_2_n10 ), .ZN(Red_ShiftRowsOutput[38]) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U7  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_2_n9 ), .A2(StateRegOutput[51]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_2_n10 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U6  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_2_n8 ), .A2(StateRegOutput[50]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_2_n9 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U5  ( .A1(StateRegOutput[48]), 
        .A2(StateRegOutput[49]), .ZN(\Red_SubCellInst_LFInst_12_LFInst_2_n8 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U4  ( .A1(StateRegOutput[49]), 
        .A2(\Red_SubCellInst_LFInst_12_LFInst_2_n7 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_2_n11 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U3  ( .A(StateRegOutput[50]), 
        .B(StateRegOutput[48]), .ZN(\Red_SubCellInst_LFInst_12_LFInst_2_n7 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U7  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_0_n8 ), .A2(
        \Red_SubCellInst_LFInst_13_LFInst_0_n7 ), .ZN(Red_ShiftRowsOutput[39])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U6  ( .A1(StateRegOutput[54]), 
        .A2(StateRegOutput[55]), .ZN(\Red_SubCellInst_LFInst_13_LFInst_0_n7 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U5  ( .A1(StateRegOutput[52]), 
        .A2(\Red_SubCellInst_LFInst_13_LFInst_0_n6 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_0_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U4  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_0_n5 ), .A2(StateRegOutput[54]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_0_n6 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U3  ( .A(StateRegOutput[53]), 
        .B(StateRegOutput[55]), .ZN(\Red_SubCellInst_LFInst_13_LFInst_0_n5 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_1_U5  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_1_n4 ), .A2(
        \Red_SubCellInst_LFInst_13_LFInst_1_n3 ), .ZN(Red_ShiftRowsOutput[40])
         );
  OR2_X1 \Red_SubCellInst_LFInst_13_LFInst_1_U4  ( .A1(StateRegOutput[55]), 
        .A2(StateRegOutput[54]), .ZN(\Red_SubCellInst_LFInst_13_LFInst_1_n3 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_1_U3  ( .A1(StateRegOutput[53]), 
        .A2(StateRegOutput[55]), .ZN(\Red_SubCellInst_LFInst_13_LFInst_1_n4 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U8  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_2_n11 ), .A2(
        \Red_SubCellInst_LFInst_13_LFInst_2_n10 ), .ZN(Red_ShiftRowsOutput[41]) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U7  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_2_n9 ), .A2(StateRegOutput[55]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_2_n10 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U6  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_2_n8 ), .A2(StateRegOutput[54]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_2_n9 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U5  ( .A1(StateRegOutput[52]), 
        .A2(StateRegOutput[53]), .ZN(\Red_SubCellInst_LFInst_13_LFInst_2_n8 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U4  ( .A1(StateRegOutput[53]), 
        .A2(\Red_SubCellInst_LFInst_13_LFInst_2_n7 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_2_n11 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U3  ( .A(StateRegOutput[54]), 
        .B(StateRegOutput[52]), .ZN(\Red_SubCellInst_LFInst_13_LFInst_2_n7 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U7  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_0_n8 ), .A2(
        \Red_SubCellInst_LFInst_14_LFInst_0_n7 ), .ZN(Red_ShiftRowsOutput[42])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U6  ( .A1(AddConstOutput[26]), 
        .A2(AddConstOutput[27]), .ZN(\Red_SubCellInst_LFInst_14_LFInst_0_n7 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U5  ( .A1(AddConstOutput[24]), 
        .A2(\Red_SubCellInst_LFInst_14_LFInst_0_n6 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_0_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U4  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_0_n5 ), .A2(AddConstOutput[26]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_0_n6 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U3  ( .A(AddConstOutput[25]), 
        .B(AddConstOutput[27]), .ZN(\Red_SubCellInst_LFInst_14_LFInst_0_n5 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_1_U5  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_1_n4 ), .A2(
        \Red_SubCellInst_LFInst_14_LFInst_1_n3 ), .ZN(Red_ShiftRowsOutput[43])
         );
  OR2_X1 \Red_SubCellInst_LFInst_14_LFInst_1_U4  ( .A1(AddConstOutput[27]), 
        .A2(AddConstOutput[26]), .ZN(\Red_SubCellInst_LFInst_14_LFInst_1_n3 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_1_U3  ( .A1(AddConstOutput[25]), 
        .A2(AddConstOutput[27]), .ZN(\Red_SubCellInst_LFInst_14_LFInst_1_n4 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U8  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_2_n11 ), .A2(
        \Red_SubCellInst_LFInst_14_LFInst_2_n10 ), .ZN(Red_ShiftRowsOutput[44]) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U7  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_2_n9 ), .A2(AddConstOutput[27]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_2_n10 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U6  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_2_n8 ), .A2(AddConstOutput[26]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_2_n9 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U5  ( .A1(AddConstOutput[24]), 
        .A2(AddConstOutput[25]), .ZN(\Red_SubCellInst_LFInst_14_LFInst_2_n8 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U4  ( .A1(AddConstOutput[25]), 
        .A2(\Red_SubCellInst_LFInst_14_LFInst_2_n7 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_2_n11 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U3  ( .A(AddConstOutput[26]), 
        .B(AddConstOutput[24]), .ZN(\Red_SubCellInst_LFInst_14_LFInst_2_n7 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U7  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_0_n8 ), .A2(
        \Red_SubCellInst_LFInst_15_LFInst_0_n7 ), .ZN(Red_ShiftRowsOutput[45])
         );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U6  ( .A1(AddConstOutput[30]), 
        .A2(AddConstOutput[31]), .ZN(\Red_SubCellInst_LFInst_15_LFInst_0_n7 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U5  ( .A1(AddConstOutput[28]), 
        .A2(\Red_SubCellInst_LFInst_15_LFInst_0_n6 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_0_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U4  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_0_n5 ), .A2(AddConstOutput[30]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_0_n6 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U3  ( .A(AddConstOutput[29]), 
        .B(AddConstOutput[31]), .ZN(\Red_SubCellInst_LFInst_15_LFInst_0_n5 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_1_U5  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_1_n4 ), .A2(
        \Red_SubCellInst_LFInst_15_LFInst_1_n3 ), .ZN(Red_ShiftRowsOutput[46])
         );
  OR2_X1 \Red_SubCellInst_LFInst_15_LFInst_1_U4  ( .A1(AddConstOutput[31]), 
        .A2(AddConstOutput[30]), .ZN(\Red_SubCellInst_LFInst_15_LFInst_1_n3 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_1_U3  ( .A1(AddConstOutput[29]), 
        .A2(AddConstOutput[31]), .ZN(\Red_SubCellInst_LFInst_15_LFInst_1_n4 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U8  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_2_n11 ), .A2(
        \Red_SubCellInst_LFInst_15_LFInst_2_n10 ), .ZN(Red_ShiftRowsOutput[47]) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U7  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_2_n9 ), .A2(AddConstOutput[31]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_2_n10 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U6  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_2_n8 ), .A2(AddConstOutput[30]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_2_n9 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U5  ( .A1(AddConstOutput[28]), 
        .A2(AddConstOutput[29]), .ZN(\Red_SubCellInst_LFInst_15_LFInst_2_n8 )
         );
  OR2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U4  ( .A1(AddConstOutput[29]), 
        .A2(\Red_SubCellInst_LFInst_15_LFInst_2_n7 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_2_n11 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U3  ( .A(AddConstOutput[30]), 
        .B(AddConstOutput[28]), .ZN(\Red_SubCellInst_LFInst_15_LFInst_2_n7 )
         );
  XOR2_X1 \Red_MCInst_MC0_v0_2Inst_0_U3  ( .A(\MCInst_MC0_v0_3 [3]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\Red_MCInst_MC0_v0_2 [0]) );
  XOR2_X1 \Red_MCInst_MC0_v0_3Inst_0_U3  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(
        \Red_MCInst_MC0_v0_2 [2]), .Z(\Red_MCInst_MC0_v0_3 [0]) );
  XNOR2_X1 \Red_MCInst_MC0_v1_0Inst_0_U4  ( .A(\Red_MCInst_MC0_v1_0Inst_0_n2 ), 
        .B(\Red_MCInst_MC0_v1_2 [1]), .ZN(\Red_MCInst_MC0_v1_0 [0]) );
  XNOR2_X1 \Red_MCInst_MC0_v1_0Inst_0_U3  ( .A(\MCInst_MC0_v1_3 [3]), .B(
        \MCInst_MC0_v1_0 [0]), .ZN(\Red_MCInst_MC0_v1_0Inst_0_n2 ) );
  XOR2_X1 \Red_MCInst_MC0_v1_2Inst_0_U3  ( .A(\Red_MCInst_MC0_v1_2 [1]), .B(
        \Red_MCInst_MC0_v1_1 [2]), .Z(\Red_MCInst_MC0_v1_2 [0]) );
  XOR2_X1 \Red_MCInst_MC0_v1_3Inst_0_U3  ( .A(\MCInst_MC0_v1_0 [0]), .B(
        \Red_MCInst_MC0_v1_2 [1]), .Z(\Red_MCInst_MC0_v1_3 [0]) );
  XOR2_X1 \Red_MCInst_MC0_v2_0Inst_0_U3  ( .A(\Red_MCInst_MC0_v2_1 [1]), .B(
        \MCInst_MC0_v2_0 [2]), .Z(\Red_MCInst_MC0_v2_0 [0]) );
  XOR2_X1 \Red_MCInst_MC0_v2_1Inst_0_U3  ( .A(\MCInst_MC0_v2_0 [2]), .B(
        \MCInst_MC0_v2_0 [3]), .Z(\Red_MCInst_MC0_v2_1 [0]) );
  XNOR2_X1 \Red_MCInst_MC0_v2_2Inst_0_U4  ( .A(\Red_MCInst_MC0_v2_2Inst_0_n2 ), 
        .B(\MCInst_MC0_v2_0 [2]), .ZN(\Red_MCInst_MC0_v2_2 [0]) );
  XNOR2_X1 \Red_MCInst_MC0_v2_2Inst_0_U3  ( .A(\Red_MCInst_MC0_v2_2 [1]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\Red_MCInst_MC0_v2_2Inst_0_n2 ) );
  XNOR2_X1 \Red_MCInst_MC0_v2_3Inst_0_U4  ( .A(\Red_MCInst_MC0_v2_3Inst_0_n2 ), 
        .B(\MCInst_MC0_v2_0 [3]), .ZN(\Red_MCInst_MC0_v2_3 [0]) );
  XNOR2_X1 \Red_MCInst_MC0_v2_3Inst_0_U3  ( .A(\Red_MCInst_MC0_v2_2 [1]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\Red_MCInst_MC0_v2_3Inst_0_n2 ) );
  XOR2_X1 \Red_MCInst_MC0_v3_0Inst_0_U3  ( .A(\MCInst_MC0_v3_2 [3]), .B(
        \Red_MCInst_MC0_v3_3 [2]), .Z(\Red_MCInst_MC0_v3_0 [0]) );
  XNOR2_X1 \Red_MCInst_MC0_v3_2Inst_0_U5  ( .A(\Red_MCInst_MC0_v3_2Inst_0_n4 ), 
        .B(\Red_MCInst_MC0_v3_2Inst_0_n3 ), .ZN(\Red_MCInst_MC0_v3_2 [0]) );
  XNOR2_X1 \Red_MCInst_MC0_v3_2Inst_0_U4  ( .A(\Red_MCInst_MC0_v3_3 [2]), .B(
        \MCInst_MC0_v3_2 [3]), .ZN(\Red_MCInst_MC0_v3_2Inst_0_n3 ) );
  XOR2_X1 \Red_MCInst_MC0_v3_2Inst_0_U3  ( .A(\MCInst_MC0_v3_0 [3]), .B(
        \Red_MCInst_MC0_v3_1 [2]), .Z(\Red_MCInst_MC0_v3_2Inst_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_v3_3Inst_0_U3  ( .A(\MCInst_MC0_v3_0 [3]), .B(
        \Red_MCInst_MC0_v3_1 [2]), .Z(\Red_MCInst_MC0_v3_3 [0]) );
  XOR2_X1 \Red_MCInst_MC0_v0_0Inst_1_U3  ( .A(\Red_MCInst_MC0_v0_2 [2]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\Red_MCInst_MC0_v0_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC0_v0_1Inst_1_U4  ( .A(\Red_MCInst_MC0_v0_1Inst_1_n2 ), 
        .B(\MCInst_MC0_v0_3 [3]), .ZN(\Red_MCInst_MC0_v0_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC0_v0_1Inst_1_U3  ( .A(\Red_MCInst_MC0_v0_1 [0]), .B(
        \Red_MCInst_MC0_v0_0 [0]), .ZN(\Red_MCInst_MC0_v0_1Inst_1_n2 ) );
  XOR2_X1 \Red_MCInst_MC0_v0_2Inst_1_U3  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(
        \Red_MCInst_MC0_v0_2 [2]), .Z(\Red_MCInst_MC0_v0_2 [1]) );
  XOR2_X1 \Red_MCInst_MC0_v0_3Inst_1_U3  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(
        \MCInst_MC0_v0_3 [3]), .Z(\Red_MCInst_MC0_v0_3 [1]) );
  XNOR2_X1 \Red_MCInst_MC0_v1_0Inst_1_U4  ( .A(\Red_MCInst_MC0_v1_0Inst_1_n2 ), 
        .B(\Red_MCInst_MC0_v1_2 [1]), .ZN(\Red_MCInst_MC0_v1_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC0_v1_0Inst_1_U3  ( .A(\Red_MCInst_MC0_v1_1 [2]), .B(
        \MCInst_MC0_v1_0 [0]), .ZN(\Red_MCInst_MC0_v1_0Inst_1_n2 ) );
  XNOR2_X1 \Red_MCInst_MC0_v1_1Inst_1_U5  ( .A(\Red_MCInst_MC0_v1_1Inst_1_n4 ), 
        .B(\Red_MCInst_MC0_v1_1Inst_1_n3 ), .ZN(\Red_MCInst_MC0_v1_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC0_v1_1Inst_1_U4  ( .A(\Red_MCInst_MC0_v1_2 [1]), .B(
        \MCInst_MC0_v1_0 [0]), .ZN(\Red_MCInst_MC0_v1_1Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_MC0_v1_1Inst_1_U3  ( .A(\MCInst_MC0_v1_3 [3]), .B(
        \Red_MCInst_MC0_v1_1 [2]), .Z(\Red_MCInst_MC0_v1_1Inst_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_v1_3Inst_1_U3  ( .A(\MCInst_MC0_v1_0 [0]), .B(
        \MCInst_MC0_v1_3 [3]), .Z(\Red_MCInst_MC0_v1_3 [1]) );
  XOR2_X1 \Red_MCInst_MC0_v2_0Inst_1_U3  ( .A(\Red_MCInst_MC0_v2_1 [1]), .B(
        \MCInst_MC0_v2_0 [3]), .Z(\Red_MCInst_MC0_v2_0 [1]) );
  XOR2_X1 \Red_MCInst_MC0_v2_3Inst_1_U3  ( .A(\Red_MCInst_MC0_v2_1 [1]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\Red_MCInst_MC0_v2_3 [1]) );
  XOR2_X1 \Red_MCInst_MC0_v3_0Inst_1_U3  ( .A(\MCInst_MC0_v3_2 [3]), .B(
        \MCInst_MC0_v3_0 [3]), .Z(\Red_MCInst_MC0_v3_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC0_v3_1Inst_1_U5  ( .A(\Red_MCInst_MC0_v3_1Inst_1_n4 ), 
        .B(\Red_MCInst_MC0_v3_1Inst_1_n3 ), .ZN(\Red_MCInst_MC0_v3_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC0_v3_1Inst_1_U4  ( .A(\Red_MCInst_MC0_v3_3 [2]), .B(
        \MCInst_MC0_v3_2 [3]), .ZN(\Red_MCInst_MC0_v3_1Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_MC0_v3_1Inst_1_U3  ( .A(\MCInst_MC0_v3_0 [3]), .B(
        \Red_MCInst_MC0_v3_1 [2]), .Z(\Red_MCInst_MC0_v3_1Inst_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_v3_2Inst_1_U3  ( .A(\Red_MCInst_MC0_v3_3 [2]), .B(
        \MCInst_MC0_v3_0 [3]), .Z(\Red_MCInst_MC0_v3_2 [1]) );
  XOR2_X1 \Red_MCInst_MC0_v3_3Inst_1_U3  ( .A(\MCInst_MC0_v3_2 [3]), .B(
        \Red_MCInst_MC0_v3_3 [2]), .Z(\Red_MCInst_MC0_v3_3 [1]) );
  XNOR2_X1 \Red_MCInst_MC0_v0_0Inst_2_U4  ( .A(\Red_MCInst_MC0_v0_0Inst_2_n2 ), 
        .B(\Red_MCInst_MC0_v0_2 [2]), .ZN(\Red_MCInst_MC0_v0_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v0_0Inst_2_U3  ( .A(\MCInst_MC0_v0_3 [3]), .B(
        \Red_MCInst_MC0_v0_0 [0]), .ZN(\Red_MCInst_MC0_v0_0Inst_2_n2 ) );
  XOR2_X1 \Red_MCInst_MC0_v0_1Inst_2_U3  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(
        \Red_MCInst_MC0_v0_2 [2]), .Z(\Red_MCInst_MC0_v0_1 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v0_3Inst_2_U5  ( .A(\Red_MCInst_MC0_v0_3Inst_2_n4 ), 
        .B(\Red_MCInst_MC0_v0_3Inst_2_n3 ), .ZN(\Red_MCInst_MC0_v0_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v0_3Inst_2_U4  ( .A(\Red_MCInst_MC0_v0_2 [2]), .B(
        \Red_MCInst_MC0_v0_0 [0]), .ZN(\Red_MCInst_MC0_v0_3Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC0_v0_3Inst_2_U3  ( .A(\MCInst_MC0_v0_3 [3]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\Red_MCInst_MC0_v0_3Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC0_v1_0Inst_2_U4  ( .A(\Red_MCInst_MC0_v1_0Inst_2_n2 ), 
        .B(\MCInst_MC0_v1_3 [3]), .ZN(\Red_MCInst_MC0_v1_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v1_0Inst_2_U3  ( .A(\Red_MCInst_MC0_v1_1 [2]), .B(
        \Red_MCInst_MC0_v1_2 [1]), .ZN(\Red_MCInst_MC0_v1_0Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC0_v1_2Inst_2_U4  ( .A(\Red_MCInst_MC0_v1_2Inst_2_n2 ), 
        .B(\Red_MCInst_MC0_v1_2 [1]), .ZN(\Red_MCInst_MC0_v1_2 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v1_2Inst_2_U3  ( .A(\Red_MCInst_MC0_v1_1 [2]), .B(
        \MCInst_MC0_v1_0 [0]), .ZN(\Red_MCInst_MC0_v1_2Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC0_v1_3Inst_2_U5  ( .A(\Red_MCInst_MC0_v1_3Inst_2_n4 ), 
        .B(\Red_MCInst_MC0_v1_3Inst_2_n3 ), .ZN(\Red_MCInst_MC0_v1_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v1_3Inst_2_U4  ( .A(\Red_MCInst_MC0_v1_2 [1]), .B(
        \MCInst_MC0_v1_0 [0]), .ZN(\Red_MCInst_MC0_v1_3Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC0_v1_3Inst_2_U3  ( .A(\MCInst_MC0_v1_3 [3]), .B(
        \Red_MCInst_MC0_v1_1 [2]), .Z(\Red_MCInst_MC0_v1_3Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC0_v2_0Inst_2_U5  ( .A(\Red_MCInst_MC0_v2_0Inst_2_n4 ), 
        .B(\Red_MCInst_MC0_v2_0Inst_2_n3 ), .ZN(\Red_MCInst_MC0_v2_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v2_0Inst_2_U4  ( .A(\MCInst_MC0_v2_0 [2]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\Red_MCInst_MC0_v2_0Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC0_v2_0Inst_2_U3  ( .A(\MCInst_MC0_v2_0 [3]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\Red_MCInst_MC0_v2_0Inst_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_v2_1Inst_2_U3  ( .A(\Red_MCInst_MC0_v2_1 [1]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\Red_MCInst_MC0_v2_1 [2]) );
  XOR2_X1 \Red_MCInst_MC0_v2_2Inst_2_U3  ( .A(\MCInst_MC0_v2_0 [3]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\Red_MCInst_MC0_v2_2 [2]) );
  XOR2_X1 \Red_MCInst_MC0_v2_3Inst_2_U3  ( .A(\Red_MCInst_MC0_v2_1 [1]), .B(
        \MCInst_MC0_v2_0 [3]), .Z(\Red_MCInst_MC0_v2_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v3_0Inst_2_U5  ( .A(\Red_MCInst_MC0_v3_0Inst_2_n4 ), 
        .B(\Red_MCInst_MC0_v3_0Inst_2_n3 ), .ZN(\Red_MCInst_MC0_v3_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v3_0Inst_2_U4  ( .A(\Red_MCInst_MC0_v3_3 [2]), .B(
        \MCInst_MC0_v3_2 [3]), .ZN(\Red_MCInst_MC0_v3_0Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC0_v3_0Inst_2_U3  ( .A(\MCInst_MC0_v3_0 [3]), .B(
        \Red_MCInst_MC0_v3_1 [2]), .Z(\Red_MCInst_MC0_v3_0Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC0_v3_2Inst_2_U4  ( .A(\Red_MCInst_MC0_v3_2Inst_2_n2 ), 
        .B(\MCInst_MC0_v3_0 [3]), .ZN(\Red_MCInst_MC0_v3_2 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v3_2Inst_2_U3  ( .A(\Red_MCInst_MC0_v3_1 [2]), .B(
        \MCInst_MC0_v3_2 [3]), .ZN(\Red_MCInst_MC0_v3_2Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC0_r0Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC0_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[45]) );
  XNOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC0_v3_0 [0]), .B(\Red_MCInst_MC0_v2_0 [0]), .ZN(
        \Red_MCInst_MC0_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(\Red_MCInst_MC0_v1_0 [0]), .Z(\Red_MCInst_MC0_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC0_r0Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC0_r0Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[46]) );
  XNOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC0_v3_0 [1]), .B(\Red_MCInst_MC0_v2_0 [1]), .ZN(
        \Red_MCInst_MC0_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC0_v0_0 [1]), .B(\Red_MCInst_MC0_v1_0 [1]), .Z(\Red_MCInst_MC0_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC0_r0Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC0_r0Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[47]) );
  XNOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC0_v3_0 [2]), .B(\Red_MCInst_MC0_v2_0 [2]), .ZN(
        \Red_MCInst_MC0_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC0_v0_0 [2]), .B(\Red_MCInst_MC0_v1_0 [2]), .Z(\Red_MCInst_MC0_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC0_r1Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC0_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[33]) );
  XNOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC0_v3_3 [2]), .B(\Red_MCInst_MC0_v2_1 [0]), .ZN(
        \Red_MCInst_MC0_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC0_v0_1 [0]), .B(\Red_MCInst_MC0_v1_2 [1]), .Z(\Red_MCInst_MC0_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC0_r1Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC0_r1Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[34]) );
  XNOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC0_v3_1 [1]), .B(\Red_MCInst_MC0_v2_1 [1]), .ZN(
        \Red_MCInst_MC0_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC0_v0_1 [1]), .B(\Red_MCInst_MC0_v1_1 [1]), .Z(\Red_MCInst_MC0_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC0_r1Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC0_r1Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[35]) );
  XNOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC0_v3_1 [2]), .B(\Red_MCInst_MC0_v2_1 [2]), .ZN(
        \Red_MCInst_MC0_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC0_v0_1 [2]), .B(\Red_MCInst_MC0_v1_1 [2]), .Z(\Red_MCInst_MC0_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC0_r2Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC0_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[21]) );
  XNOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC0_v3_2 [0]), .B(\Red_MCInst_MC0_v2_2 [0]), .ZN(
        \Red_MCInst_MC0_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC0_v0_2 [0]), .B(\Red_MCInst_MC0_v1_2 [0]), .Z(\Red_MCInst_MC0_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC0_r2Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC0_r2Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[22]) );
  XNOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC0_v3_2 [1]), .B(\Red_MCInst_MC0_v2_2 [1]), .ZN(
        \Red_MCInst_MC0_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC0_v0_2 [1]), .B(\Red_MCInst_MC0_v1_2 [1]), .Z(\Red_MCInst_MC0_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC0_r2Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC0_r2Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[23]) );
  XNOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC0_v3_2 [2]), .B(\Red_MCInst_MC0_v2_2 [2]), .ZN(
        \Red_MCInst_MC0_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC0_v0_2 [2]), .B(\Red_MCInst_MC0_v1_2 [2]), .Z(\Red_MCInst_MC0_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC0_r3Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC0_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[9]) );
  XNOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC0_v3_3 [0]), .B(\Red_MCInst_MC0_v2_3 [0]), .ZN(
        \Red_MCInst_MC0_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC0_v0_3 [0]), .B(\Red_MCInst_MC0_v1_3 [0]), .Z(\Red_MCInst_MC0_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC0_r3Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC0_r3Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[10]) );
  XNOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC0_v3_3 [1]), .B(\Red_MCInst_MC0_v2_3 [1]), .ZN(
        \Red_MCInst_MC0_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC0_v0_3 [1]), .B(\Red_MCInst_MC0_v1_3 [1]), .Z(\Red_MCInst_MC0_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC0_r3Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC0_r3Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[11]) );
  XNOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC0_v3_3 [2]), .B(\Red_MCInst_MC0_v2_3 [2]), .ZN(
        \Red_MCInst_MC0_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC0_v0_3 [2]), .B(\Red_MCInst_MC0_v1_3 [2]), .Z(\Red_MCInst_MC0_r3Inst_XORInst_0_2_n5 ) );
  XOR2_X1 \Red_MCInst_MC1_v0_2Inst_0_U3  ( .A(\MCInst_MC1_v0_3 [3]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\Red_MCInst_MC1_v0_2 [0]) );
  XOR2_X1 \Red_MCInst_MC1_v0_3Inst_0_U3  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(
        \Red_MCInst_MC1_v0_2 [2]), .Z(\Red_MCInst_MC1_v0_3 [0]) );
  XNOR2_X1 \Red_MCInst_MC1_v1_0Inst_0_U4  ( .A(\Red_MCInst_MC1_v1_0Inst_0_n2 ), 
        .B(\Red_MCInst_MC1_v1_2 [1]), .ZN(\Red_MCInst_MC1_v1_0 [0]) );
  XNOR2_X1 \Red_MCInst_MC1_v1_0Inst_0_U3  ( .A(\MCInst_MC1_v1_3 [3]), .B(
        \MCInst_MC1_v1_0 [0]), .ZN(\Red_MCInst_MC1_v1_0Inst_0_n2 ) );
  XOR2_X1 \Red_MCInst_MC1_v1_2Inst_0_U3  ( .A(\Red_MCInst_MC1_v1_2 [1]), .B(
        \Red_MCInst_MC1_v1_1 [2]), .Z(\Red_MCInst_MC1_v1_2 [0]) );
  XOR2_X1 \Red_MCInst_MC1_v1_3Inst_0_U3  ( .A(\MCInst_MC1_v1_0 [0]), .B(
        \Red_MCInst_MC1_v1_2 [1]), .Z(\Red_MCInst_MC1_v1_3 [0]) );
  XOR2_X1 \Red_MCInst_MC1_v2_0Inst_0_U3  ( .A(\Red_MCInst_MC1_v2_1 [1]), .B(
        \MCInst_MC1_v2_0 [2]), .Z(\Red_MCInst_MC1_v2_0 [0]) );
  XOR2_X1 \Red_MCInst_MC1_v2_1Inst_0_U3  ( .A(\MCInst_MC1_v2_0 [2]), .B(
        \MCInst_MC1_v2_0 [3]), .Z(\Red_MCInst_MC1_v2_1 [0]) );
  XNOR2_X1 \Red_MCInst_MC1_v2_2Inst_0_U4  ( .A(\Red_MCInst_MC1_v2_2Inst_0_n2 ), 
        .B(\MCInst_MC1_v2_0 [2]), .ZN(\Red_MCInst_MC1_v2_2 [0]) );
  XNOR2_X1 \Red_MCInst_MC1_v2_2Inst_0_U3  ( .A(\Red_MCInst_MC1_v2_2 [1]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\Red_MCInst_MC1_v2_2Inst_0_n2 ) );
  XNOR2_X1 \Red_MCInst_MC1_v2_3Inst_0_U4  ( .A(\Red_MCInst_MC1_v2_3Inst_0_n2 ), 
        .B(\MCInst_MC1_v2_0 [3]), .ZN(\Red_MCInst_MC1_v2_3 [0]) );
  XNOR2_X1 \Red_MCInst_MC1_v2_3Inst_0_U3  ( .A(\Red_MCInst_MC1_v2_2 [1]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\Red_MCInst_MC1_v2_3Inst_0_n2 ) );
  XOR2_X1 \Red_MCInst_MC1_v3_0Inst_0_U3  ( .A(\MCInst_MC1_v3_2 [3]), .B(
        \Red_MCInst_MC1_v3_3 [2]), .Z(\Red_MCInst_MC1_v3_0 [0]) );
  XNOR2_X1 \Red_MCInst_MC1_v3_2Inst_0_U5  ( .A(\Red_MCInst_MC1_v3_2Inst_0_n4 ), 
        .B(\Red_MCInst_MC1_v3_2Inst_0_n3 ), .ZN(\Red_MCInst_MC1_v3_2 [0]) );
  XNOR2_X1 \Red_MCInst_MC1_v3_2Inst_0_U4  ( .A(\Red_MCInst_MC1_v3_3 [2]), .B(
        \MCInst_MC1_v3_2 [3]), .ZN(\Red_MCInst_MC1_v3_2Inst_0_n3 ) );
  XOR2_X1 \Red_MCInst_MC1_v3_2Inst_0_U3  ( .A(\MCInst_MC1_v3_0 [3]), .B(
        \Red_MCInst_MC1_v3_1 [2]), .Z(\Red_MCInst_MC1_v3_2Inst_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_v3_3Inst_0_U3  ( .A(\MCInst_MC1_v3_0 [3]), .B(
        \Red_MCInst_MC1_v3_1 [2]), .Z(\Red_MCInst_MC1_v3_3 [0]) );
  XOR2_X1 \Red_MCInst_MC1_v0_0Inst_1_U3  ( .A(\Red_MCInst_MC1_v0_2 [2]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\Red_MCInst_MC1_v0_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC1_v0_1Inst_1_U4  ( .A(\Red_MCInst_MC1_v0_1Inst_1_n2 ), 
        .B(\MCInst_MC1_v0_3 [3]), .ZN(\Red_MCInst_MC1_v0_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC1_v0_1Inst_1_U3  ( .A(\Red_MCInst_MC1_v0_1 [0]), .B(
        \Red_MCInst_MC1_v0_0 [0]), .ZN(\Red_MCInst_MC1_v0_1Inst_1_n2 ) );
  XOR2_X1 \Red_MCInst_MC1_v0_2Inst_1_U3  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(
        \Red_MCInst_MC1_v0_2 [2]), .Z(\Red_MCInst_MC1_v0_2 [1]) );
  XOR2_X1 \Red_MCInst_MC1_v0_3Inst_1_U3  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(
        \MCInst_MC1_v0_3 [3]), .Z(\Red_MCInst_MC1_v0_3 [1]) );
  XNOR2_X1 \Red_MCInst_MC1_v1_0Inst_1_U4  ( .A(\Red_MCInst_MC1_v1_0Inst_1_n2 ), 
        .B(\Red_MCInst_MC1_v1_2 [1]), .ZN(\Red_MCInst_MC1_v1_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC1_v1_0Inst_1_U3  ( .A(\Red_MCInst_MC1_v1_1 [2]), .B(
        \MCInst_MC1_v1_0 [0]), .ZN(\Red_MCInst_MC1_v1_0Inst_1_n2 ) );
  XNOR2_X1 \Red_MCInst_MC1_v1_1Inst_1_U5  ( .A(\Red_MCInst_MC1_v1_1Inst_1_n4 ), 
        .B(\Red_MCInst_MC1_v1_1Inst_1_n3 ), .ZN(\Red_MCInst_MC1_v1_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC1_v1_1Inst_1_U4  ( .A(\Red_MCInst_MC1_v1_2 [1]), .B(
        \MCInst_MC1_v1_0 [0]), .ZN(\Red_MCInst_MC1_v1_1Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_MC1_v1_1Inst_1_U3  ( .A(\MCInst_MC1_v1_3 [3]), .B(
        \Red_MCInst_MC1_v1_1 [2]), .Z(\Red_MCInst_MC1_v1_1Inst_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_v1_3Inst_1_U3  ( .A(\MCInst_MC1_v1_0 [0]), .B(
        \MCInst_MC1_v1_3 [3]), .Z(\Red_MCInst_MC1_v1_3 [1]) );
  XOR2_X1 \Red_MCInst_MC1_v2_0Inst_1_U3  ( .A(\Red_MCInst_MC1_v2_1 [1]), .B(
        \MCInst_MC1_v2_0 [3]), .Z(\Red_MCInst_MC1_v2_0 [1]) );
  XOR2_X1 \Red_MCInst_MC1_v2_3Inst_1_U3  ( .A(\Red_MCInst_MC1_v2_1 [1]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\Red_MCInst_MC1_v2_3 [1]) );
  XOR2_X1 \Red_MCInst_MC1_v3_0Inst_1_U3  ( .A(\MCInst_MC1_v3_2 [3]), .B(
        \MCInst_MC1_v3_0 [3]), .Z(\Red_MCInst_MC1_v3_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC1_v3_1Inst_1_U5  ( .A(\Red_MCInst_MC1_v3_1Inst_1_n4 ), 
        .B(\Red_MCInst_MC1_v3_1Inst_1_n3 ), .ZN(\Red_MCInst_MC1_v3_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC1_v3_1Inst_1_U4  ( .A(\Red_MCInst_MC1_v3_3 [2]), .B(
        \MCInst_MC1_v3_2 [3]), .ZN(\Red_MCInst_MC1_v3_1Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_MC1_v3_1Inst_1_U3  ( .A(\MCInst_MC1_v3_0 [3]), .B(
        \Red_MCInst_MC1_v3_1 [2]), .Z(\Red_MCInst_MC1_v3_1Inst_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_v3_2Inst_1_U3  ( .A(\Red_MCInst_MC1_v3_3 [2]), .B(
        \MCInst_MC1_v3_0 [3]), .Z(\Red_MCInst_MC1_v3_2 [1]) );
  XOR2_X1 \Red_MCInst_MC1_v3_3Inst_1_U3  ( .A(\MCInst_MC1_v3_2 [3]), .B(
        \Red_MCInst_MC1_v3_3 [2]), .Z(\Red_MCInst_MC1_v3_3 [1]) );
  XNOR2_X1 \Red_MCInst_MC1_v0_0Inst_2_U4  ( .A(\Red_MCInst_MC1_v0_0Inst_2_n2 ), 
        .B(\Red_MCInst_MC1_v0_2 [2]), .ZN(\Red_MCInst_MC1_v0_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v0_0Inst_2_U3  ( .A(\MCInst_MC1_v0_3 [3]), .B(
        \Red_MCInst_MC1_v0_0 [0]), .ZN(\Red_MCInst_MC1_v0_0Inst_2_n2 ) );
  XOR2_X1 \Red_MCInst_MC1_v0_1Inst_2_U3  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(
        \Red_MCInst_MC1_v0_2 [2]), .Z(\Red_MCInst_MC1_v0_1 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v0_3Inst_2_U5  ( .A(\Red_MCInst_MC1_v0_3Inst_2_n4 ), 
        .B(\Red_MCInst_MC1_v0_3Inst_2_n3 ), .ZN(\Red_MCInst_MC1_v0_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v0_3Inst_2_U4  ( .A(\Red_MCInst_MC1_v0_2 [2]), .B(
        \Red_MCInst_MC1_v0_0 [0]), .ZN(\Red_MCInst_MC1_v0_3Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC1_v0_3Inst_2_U3  ( .A(\MCInst_MC1_v0_3 [3]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\Red_MCInst_MC1_v0_3Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC1_v1_0Inst_2_U4  ( .A(\Red_MCInst_MC1_v1_0Inst_2_n2 ), 
        .B(\MCInst_MC1_v1_3 [3]), .ZN(\Red_MCInst_MC1_v1_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v1_0Inst_2_U3  ( .A(\Red_MCInst_MC1_v1_1 [2]), .B(
        \Red_MCInst_MC1_v1_2 [1]), .ZN(\Red_MCInst_MC1_v1_0Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC1_v1_2Inst_2_U4  ( .A(\Red_MCInst_MC1_v1_2Inst_2_n2 ), 
        .B(\Red_MCInst_MC1_v1_2 [1]), .ZN(\Red_MCInst_MC1_v1_2 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v1_2Inst_2_U3  ( .A(\Red_MCInst_MC1_v1_1 [2]), .B(
        \MCInst_MC1_v1_0 [0]), .ZN(\Red_MCInst_MC1_v1_2Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC1_v1_3Inst_2_U5  ( .A(\Red_MCInst_MC1_v1_3Inst_2_n4 ), 
        .B(\Red_MCInst_MC1_v1_3Inst_2_n3 ), .ZN(\Red_MCInst_MC1_v1_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v1_3Inst_2_U4  ( .A(\Red_MCInst_MC1_v1_2 [1]), .B(
        \MCInst_MC1_v1_0 [0]), .ZN(\Red_MCInst_MC1_v1_3Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC1_v1_3Inst_2_U3  ( .A(\MCInst_MC1_v1_3 [3]), .B(
        \Red_MCInst_MC1_v1_1 [2]), .Z(\Red_MCInst_MC1_v1_3Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC1_v2_0Inst_2_U5  ( .A(\Red_MCInst_MC1_v2_0Inst_2_n4 ), 
        .B(\Red_MCInst_MC1_v2_0Inst_2_n3 ), .ZN(\Red_MCInst_MC1_v2_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v2_0Inst_2_U4  ( .A(\MCInst_MC1_v2_0 [2]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\Red_MCInst_MC1_v2_0Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC1_v2_0Inst_2_U3  ( .A(\MCInst_MC1_v2_0 [3]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\Red_MCInst_MC1_v2_0Inst_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_v2_1Inst_2_U3  ( .A(\Red_MCInst_MC1_v2_1 [1]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\Red_MCInst_MC1_v2_1 [2]) );
  XOR2_X1 \Red_MCInst_MC1_v2_2Inst_2_U3  ( .A(\MCInst_MC1_v2_0 [3]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\Red_MCInst_MC1_v2_2 [2]) );
  XOR2_X1 \Red_MCInst_MC1_v2_3Inst_2_U3  ( .A(\Red_MCInst_MC1_v2_1 [1]), .B(
        \MCInst_MC1_v2_0 [3]), .Z(\Red_MCInst_MC1_v2_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v3_0Inst_2_U5  ( .A(\Red_MCInst_MC1_v3_0Inst_2_n4 ), 
        .B(\Red_MCInst_MC1_v3_0Inst_2_n3 ), .ZN(\Red_MCInst_MC1_v3_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v3_0Inst_2_U4  ( .A(\Red_MCInst_MC1_v3_3 [2]), .B(
        \MCInst_MC1_v3_2 [3]), .ZN(\Red_MCInst_MC1_v3_0Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC1_v3_0Inst_2_U3  ( .A(\MCInst_MC1_v3_0 [3]), .B(
        \Red_MCInst_MC1_v3_1 [2]), .Z(\Red_MCInst_MC1_v3_0Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC1_v3_2Inst_2_U4  ( .A(\Red_MCInst_MC1_v3_2Inst_2_n2 ), 
        .B(\MCInst_MC1_v3_0 [3]), .ZN(\Red_MCInst_MC1_v3_2 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v3_2Inst_2_U3  ( .A(\Red_MCInst_MC1_v3_1 [2]), .B(
        \MCInst_MC1_v3_2 [3]), .ZN(\Red_MCInst_MC1_v3_2Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC1_r0Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC1_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[42]) );
  XNOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC1_v3_0 [0]), .B(\Red_MCInst_MC1_v2_0 [0]), .ZN(
        \Red_MCInst_MC1_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(\Red_MCInst_MC1_v1_0 [0]), .Z(\Red_MCInst_MC1_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC1_r0Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC1_r0Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[43]) );
  XNOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC1_v3_0 [1]), .B(\Red_MCInst_MC1_v2_0 [1]), .ZN(
        \Red_MCInst_MC1_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC1_v0_0 [1]), .B(\Red_MCInst_MC1_v1_0 [1]), .Z(\Red_MCInst_MC1_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC1_r0Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC1_r0Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[44]) );
  XNOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC1_v3_0 [2]), .B(\Red_MCInst_MC1_v2_0 [2]), .ZN(
        \Red_MCInst_MC1_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC1_v0_0 [2]), .B(\Red_MCInst_MC1_v1_0 [2]), .Z(\Red_MCInst_MC1_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC1_r1Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC1_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[30]) );
  XNOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC1_v3_3 [2]), .B(\Red_MCInst_MC1_v2_1 [0]), .ZN(
        \Red_MCInst_MC1_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC1_v0_1 [0]), .B(\Red_MCInst_MC1_v1_2 [1]), .Z(\Red_MCInst_MC1_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC1_r1Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC1_r1Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[31]) );
  XNOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC1_v3_1 [1]), .B(\Red_MCInst_MC1_v2_1 [1]), .ZN(
        \Red_MCInst_MC1_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC1_v0_1 [1]), .B(\Red_MCInst_MC1_v1_1 [1]), .Z(\Red_MCInst_MC1_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC1_r1Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC1_r1Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[32]) );
  XNOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC1_v3_1 [2]), .B(\Red_MCInst_MC1_v2_1 [2]), .ZN(
        \Red_MCInst_MC1_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC1_v0_1 [2]), .B(\Red_MCInst_MC1_v1_1 [2]), .Z(\Red_MCInst_MC1_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC1_r2Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC1_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[18]) );
  XNOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC1_v3_2 [0]), .B(\Red_MCInst_MC1_v2_2 [0]), .ZN(
        \Red_MCInst_MC1_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC1_v0_2 [0]), .B(\Red_MCInst_MC1_v1_2 [0]), .Z(\Red_MCInst_MC1_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC1_r2Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC1_r2Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[19]) );
  XNOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC1_v3_2 [1]), .B(\Red_MCInst_MC1_v2_2 [1]), .ZN(
        \Red_MCInst_MC1_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC1_v0_2 [1]), .B(\Red_MCInst_MC1_v1_2 [1]), .Z(\Red_MCInst_MC1_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC1_r2Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC1_r2Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[20]) );
  XNOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC1_v3_2 [2]), .B(\Red_MCInst_MC1_v2_2 [2]), .ZN(
        \Red_MCInst_MC1_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC1_v0_2 [2]), .B(\Red_MCInst_MC1_v1_2 [2]), .Z(\Red_MCInst_MC1_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC1_r3Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC1_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[6]) );
  XNOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC1_v3_3 [0]), .B(\Red_MCInst_MC1_v2_3 [0]), .ZN(
        \Red_MCInst_MC1_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC1_v0_3 [0]), .B(\Red_MCInst_MC1_v1_3 [0]), .Z(\Red_MCInst_MC1_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC1_r3Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC1_r3Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[7]) );
  XNOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC1_v3_3 [1]), .B(\Red_MCInst_MC1_v2_3 [1]), .ZN(
        \Red_MCInst_MC1_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC1_v0_3 [1]), .B(\Red_MCInst_MC1_v1_3 [1]), .Z(\Red_MCInst_MC1_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC1_r3Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC1_r3Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[8]) );
  XNOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC1_v3_3 [2]), .B(\Red_MCInst_MC1_v2_3 [2]), .ZN(
        \Red_MCInst_MC1_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC1_v0_3 [2]), .B(\Red_MCInst_MC1_v1_3 [2]), .Z(\Red_MCInst_MC1_r3Inst_XORInst_0_2_n5 ) );
  XOR2_X1 \Red_MCInst_MC2_v0_2Inst_0_U3  ( .A(\MCInst_MC2_v0_3 [3]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\Red_MCInst_MC2_v0_2 [0]) );
  XOR2_X1 \Red_MCInst_MC2_v0_3Inst_0_U3  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(
        \Red_MCInst_MC2_v0_2 [2]), .Z(\Red_MCInst_MC2_v0_3 [0]) );
  XNOR2_X1 \Red_MCInst_MC2_v1_0Inst_0_U4  ( .A(\Red_MCInst_MC2_v1_0Inst_0_n2 ), 
        .B(\Red_MCInst_MC2_v1_2 [1]), .ZN(\Red_MCInst_MC2_v1_0 [0]) );
  XNOR2_X1 \Red_MCInst_MC2_v1_0Inst_0_U3  ( .A(\MCInst_MC2_v1_3 [3]), .B(
        \MCInst_MC2_v1_0 [0]), .ZN(\Red_MCInst_MC2_v1_0Inst_0_n2 ) );
  XOR2_X1 \Red_MCInst_MC2_v1_2Inst_0_U3  ( .A(\Red_MCInst_MC2_v1_2 [1]), .B(
        \Red_MCInst_MC2_v1_1 [2]), .Z(\Red_MCInst_MC2_v1_2 [0]) );
  XOR2_X1 \Red_MCInst_MC2_v1_3Inst_0_U3  ( .A(\MCInst_MC2_v1_0 [0]), .B(
        \Red_MCInst_MC2_v1_2 [1]), .Z(\Red_MCInst_MC2_v1_3 [0]) );
  XOR2_X1 \Red_MCInst_MC2_v2_0Inst_0_U3  ( .A(\Red_MCInst_MC2_v2_1 [1]), .B(
        \MCInst_MC2_v2_0 [2]), .Z(\Red_MCInst_MC2_v2_0 [0]) );
  XOR2_X1 \Red_MCInst_MC2_v2_1Inst_0_U3  ( .A(\MCInst_MC2_v2_0 [2]), .B(
        \MCInst_MC2_v2_0 [3]), .Z(\Red_MCInst_MC2_v2_1 [0]) );
  XNOR2_X1 \Red_MCInst_MC2_v2_2Inst_0_U4  ( .A(\Red_MCInst_MC2_v2_2Inst_0_n2 ), 
        .B(\MCInst_MC2_v2_0 [2]), .ZN(\Red_MCInst_MC2_v2_2 [0]) );
  XNOR2_X1 \Red_MCInst_MC2_v2_2Inst_0_U3  ( .A(\Red_MCInst_MC2_v2_2 [1]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\Red_MCInst_MC2_v2_2Inst_0_n2 ) );
  XNOR2_X1 \Red_MCInst_MC2_v2_3Inst_0_U4  ( .A(\Red_MCInst_MC2_v2_3Inst_0_n2 ), 
        .B(\MCInst_MC2_v2_0 [3]), .ZN(\Red_MCInst_MC2_v2_3 [0]) );
  XNOR2_X1 \Red_MCInst_MC2_v2_3Inst_0_U3  ( .A(\Red_MCInst_MC2_v2_2 [1]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\Red_MCInst_MC2_v2_3Inst_0_n2 ) );
  XOR2_X1 \Red_MCInst_MC2_v3_0Inst_0_U3  ( .A(\MCInst_MC2_v3_2 [3]), .B(
        \Red_MCInst_MC2_v3_3 [2]), .Z(\Red_MCInst_MC2_v3_0 [0]) );
  XNOR2_X1 \Red_MCInst_MC2_v3_2Inst_0_U5  ( .A(\Red_MCInst_MC2_v3_2Inst_0_n4 ), 
        .B(\Red_MCInst_MC2_v3_2Inst_0_n3 ), .ZN(\Red_MCInst_MC2_v3_2 [0]) );
  XNOR2_X1 \Red_MCInst_MC2_v3_2Inst_0_U4  ( .A(\Red_MCInst_MC2_v3_3 [2]), .B(
        \MCInst_MC2_v3_2 [3]), .ZN(\Red_MCInst_MC2_v3_2Inst_0_n3 ) );
  XOR2_X1 \Red_MCInst_MC2_v3_2Inst_0_U3  ( .A(\MCInst_MC2_v3_0 [3]), .B(
        \Red_MCInst_MC2_v3_1 [2]), .Z(\Red_MCInst_MC2_v3_2Inst_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_v3_3Inst_0_U3  ( .A(\MCInst_MC2_v3_0 [3]), .B(
        \Red_MCInst_MC2_v3_1 [2]), .Z(\Red_MCInst_MC2_v3_3 [0]) );
  XOR2_X1 \Red_MCInst_MC2_v0_0Inst_1_U3  ( .A(\Red_MCInst_MC2_v0_2 [2]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\Red_MCInst_MC2_v0_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC2_v0_1Inst_1_U4  ( .A(\Red_MCInst_MC2_v0_1Inst_1_n2 ), 
        .B(\MCInst_MC2_v0_3 [3]), .ZN(\Red_MCInst_MC2_v0_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC2_v0_1Inst_1_U3  ( .A(\Red_MCInst_MC2_v0_1 [0]), .B(
        \Red_MCInst_MC2_v0_0 [0]), .ZN(\Red_MCInst_MC2_v0_1Inst_1_n2 ) );
  XOR2_X1 \Red_MCInst_MC2_v0_2Inst_1_U3  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(
        \Red_MCInst_MC2_v0_2 [2]), .Z(\Red_MCInst_MC2_v0_2 [1]) );
  XOR2_X1 \Red_MCInst_MC2_v0_3Inst_1_U3  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(
        \MCInst_MC2_v0_3 [3]), .Z(\Red_MCInst_MC2_v0_3 [1]) );
  XNOR2_X1 \Red_MCInst_MC2_v1_0Inst_1_U4  ( .A(\Red_MCInst_MC2_v1_0Inst_1_n2 ), 
        .B(\Red_MCInst_MC2_v1_2 [1]), .ZN(\Red_MCInst_MC2_v1_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC2_v1_0Inst_1_U3  ( .A(\Red_MCInst_MC2_v1_1 [2]), .B(
        \MCInst_MC2_v1_0 [0]), .ZN(\Red_MCInst_MC2_v1_0Inst_1_n2 ) );
  XNOR2_X1 \Red_MCInst_MC2_v1_1Inst_1_U5  ( .A(\Red_MCInst_MC2_v1_1Inst_1_n4 ), 
        .B(\Red_MCInst_MC2_v1_1Inst_1_n3 ), .ZN(\Red_MCInst_MC2_v1_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC2_v1_1Inst_1_U4  ( .A(\Red_MCInst_MC2_v1_2 [1]), .B(
        \MCInst_MC2_v1_0 [0]), .ZN(\Red_MCInst_MC2_v1_1Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_MC2_v1_1Inst_1_U3  ( .A(\MCInst_MC2_v1_3 [3]), .B(
        \Red_MCInst_MC2_v1_1 [2]), .Z(\Red_MCInst_MC2_v1_1Inst_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_v1_3Inst_1_U3  ( .A(\MCInst_MC2_v1_0 [0]), .B(
        \MCInst_MC2_v1_3 [3]), .Z(\Red_MCInst_MC2_v1_3 [1]) );
  XOR2_X1 \Red_MCInst_MC2_v2_0Inst_1_U3  ( .A(\Red_MCInst_MC2_v2_1 [1]), .B(
        \MCInst_MC2_v2_0 [3]), .Z(\Red_MCInst_MC2_v2_0 [1]) );
  XOR2_X1 \Red_MCInst_MC2_v2_3Inst_1_U3  ( .A(\Red_MCInst_MC2_v2_1 [1]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\Red_MCInst_MC2_v2_3 [1]) );
  XOR2_X1 \Red_MCInst_MC2_v3_0Inst_1_U3  ( .A(\MCInst_MC2_v3_2 [3]), .B(
        \MCInst_MC2_v3_0 [3]), .Z(\Red_MCInst_MC2_v3_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC2_v3_1Inst_1_U5  ( .A(\Red_MCInst_MC2_v3_1Inst_1_n4 ), 
        .B(\Red_MCInst_MC2_v3_1Inst_1_n3 ), .ZN(\Red_MCInst_MC2_v3_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC2_v3_1Inst_1_U4  ( .A(\Red_MCInst_MC2_v3_3 [2]), .B(
        \MCInst_MC2_v3_2 [3]), .ZN(\Red_MCInst_MC2_v3_1Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_MC2_v3_1Inst_1_U3  ( .A(\MCInst_MC2_v3_0 [3]), .B(
        \Red_MCInst_MC2_v3_1 [2]), .Z(\Red_MCInst_MC2_v3_1Inst_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_v3_2Inst_1_U3  ( .A(\Red_MCInst_MC2_v3_3 [2]), .B(
        \MCInst_MC2_v3_0 [3]), .Z(\Red_MCInst_MC2_v3_2 [1]) );
  XOR2_X1 \Red_MCInst_MC2_v3_3Inst_1_U3  ( .A(\MCInst_MC2_v3_2 [3]), .B(
        \Red_MCInst_MC2_v3_3 [2]), .Z(\Red_MCInst_MC2_v3_3 [1]) );
  XNOR2_X1 \Red_MCInst_MC2_v0_0Inst_2_U4  ( .A(\Red_MCInst_MC2_v0_0Inst_2_n2 ), 
        .B(\Red_MCInst_MC2_v0_2 [2]), .ZN(\Red_MCInst_MC2_v0_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v0_0Inst_2_U3  ( .A(\MCInst_MC2_v0_3 [3]), .B(
        \Red_MCInst_MC2_v0_0 [0]), .ZN(\Red_MCInst_MC2_v0_0Inst_2_n2 ) );
  XOR2_X1 \Red_MCInst_MC2_v0_1Inst_2_U3  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(
        \Red_MCInst_MC2_v0_2 [2]), .Z(\Red_MCInst_MC2_v0_1 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v0_3Inst_2_U5  ( .A(\Red_MCInst_MC2_v0_3Inst_2_n4 ), 
        .B(\Red_MCInst_MC2_v0_3Inst_2_n3 ), .ZN(\Red_MCInst_MC2_v0_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v0_3Inst_2_U4  ( .A(\Red_MCInst_MC2_v0_2 [2]), .B(
        \Red_MCInst_MC2_v0_0 [0]), .ZN(\Red_MCInst_MC2_v0_3Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC2_v0_3Inst_2_U3  ( .A(\MCInst_MC2_v0_3 [3]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\Red_MCInst_MC2_v0_3Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC2_v1_0Inst_2_U4  ( .A(\Red_MCInst_MC2_v1_0Inst_2_n2 ), 
        .B(\MCInst_MC2_v1_3 [3]), .ZN(\Red_MCInst_MC2_v1_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v1_0Inst_2_U3  ( .A(\Red_MCInst_MC2_v1_1 [2]), .B(
        \Red_MCInst_MC2_v1_2 [1]), .ZN(\Red_MCInst_MC2_v1_0Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC2_v1_2Inst_2_U4  ( .A(\Red_MCInst_MC2_v1_2Inst_2_n2 ), 
        .B(\Red_MCInst_MC2_v1_2 [1]), .ZN(\Red_MCInst_MC2_v1_2 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v1_2Inst_2_U3  ( .A(\Red_MCInst_MC2_v1_1 [2]), .B(
        \MCInst_MC2_v1_0 [0]), .ZN(\Red_MCInst_MC2_v1_2Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC2_v1_3Inst_2_U5  ( .A(\Red_MCInst_MC2_v1_3Inst_2_n4 ), 
        .B(\Red_MCInst_MC2_v1_3Inst_2_n3 ), .ZN(\Red_MCInst_MC2_v1_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v1_3Inst_2_U4  ( .A(\Red_MCInst_MC2_v1_2 [1]), .B(
        \MCInst_MC2_v1_0 [0]), .ZN(\Red_MCInst_MC2_v1_3Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC2_v1_3Inst_2_U3  ( .A(\MCInst_MC2_v1_3 [3]), .B(
        \Red_MCInst_MC2_v1_1 [2]), .Z(\Red_MCInst_MC2_v1_3Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC2_v2_0Inst_2_U5  ( .A(\Red_MCInst_MC2_v2_0Inst_2_n4 ), 
        .B(\Red_MCInst_MC2_v2_0Inst_2_n3 ), .ZN(\Red_MCInst_MC2_v2_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v2_0Inst_2_U4  ( .A(\MCInst_MC2_v2_0 [2]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\Red_MCInst_MC2_v2_0Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC2_v2_0Inst_2_U3  ( .A(\MCInst_MC2_v2_0 [3]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\Red_MCInst_MC2_v2_0Inst_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_v2_1Inst_2_U3  ( .A(\Red_MCInst_MC2_v2_1 [1]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\Red_MCInst_MC2_v2_1 [2]) );
  XOR2_X1 \Red_MCInst_MC2_v2_2Inst_2_U3  ( .A(\MCInst_MC2_v2_0 [3]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\Red_MCInst_MC2_v2_2 [2]) );
  XOR2_X1 \Red_MCInst_MC2_v2_3Inst_2_U3  ( .A(\Red_MCInst_MC2_v2_1 [1]), .B(
        \MCInst_MC2_v2_0 [3]), .Z(\Red_MCInst_MC2_v2_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v3_0Inst_2_U5  ( .A(\Red_MCInst_MC2_v3_0Inst_2_n4 ), 
        .B(\Red_MCInst_MC2_v3_0Inst_2_n3 ), .ZN(\Red_MCInst_MC2_v3_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v3_0Inst_2_U4  ( .A(\Red_MCInst_MC2_v3_3 [2]), .B(
        \MCInst_MC2_v3_2 [3]), .ZN(\Red_MCInst_MC2_v3_0Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC2_v3_0Inst_2_U3  ( .A(\MCInst_MC2_v3_0 [3]), .B(
        \Red_MCInst_MC2_v3_1 [2]), .Z(\Red_MCInst_MC2_v3_0Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC2_v3_2Inst_2_U4  ( .A(\Red_MCInst_MC2_v3_2Inst_2_n2 ), 
        .B(\MCInst_MC2_v3_0 [3]), .ZN(\Red_MCInst_MC2_v3_2 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v3_2Inst_2_U3  ( .A(\Red_MCInst_MC2_v3_1 [2]), .B(
        \MCInst_MC2_v3_2 [3]), .ZN(\Red_MCInst_MC2_v3_2Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC2_r0Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC2_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[39]) );
  XNOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC2_v3_0 [0]), .B(\Red_MCInst_MC2_v2_0 [0]), .ZN(
        \Red_MCInst_MC2_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(\Red_MCInst_MC2_v1_0 [0]), .Z(\Red_MCInst_MC2_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC2_r0Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC2_r0Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[40]) );
  XNOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC2_v3_0 [1]), .B(\Red_MCInst_MC2_v2_0 [1]), .ZN(
        \Red_MCInst_MC2_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC2_v0_0 [1]), .B(\Red_MCInst_MC2_v1_0 [1]), .Z(\Red_MCInst_MC2_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC2_r0Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC2_r0Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[41]) );
  XNOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC2_v3_0 [2]), .B(\Red_MCInst_MC2_v2_0 [2]), .ZN(
        \Red_MCInst_MC2_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC2_v0_0 [2]), .B(\Red_MCInst_MC2_v1_0 [2]), .Z(\Red_MCInst_MC2_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC2_r1Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC2_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[27]) );
  XNOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC2_v3_3 [2]), .B(\Red_MCInst_MC2_v2_1 [0]), .ZN(
        \Red_MCInst_MC2_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC2_v0_1 [0]), .B(\Red_MCInst_MC2_v1_2 [1]), .Z(\Red_MCInst_MC2_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC2_r1Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC2_r1Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[28]) );
  XNOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC2_v3_1 [1]), .B(\Red_MCInst_MC2_v2_1 [1]), .ZN(
        \Red_MCInst_MC2_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC2_v0_1 [1]), .B(\Red_MCInst_MC2_v1_1 [1]), .Z(\Red_MCInst_MC2_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC2_r1Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC2_r1Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[29]) );
  XNOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC2_v3_1 [2]), .B(\Red_MCInst_MC2_v2_1 [2]), .ZN(
        \Red_MCInst_MC2_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC2_v0_1 [2]), .B(\Red_MCInst_MC2_v1_1 [2]), .Z(\Red_MCInst_MC2_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC2_r2Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC2_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[15]) );
  XNOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC2_v3_2 [0]), .B(\Red_MCInst_MC2_v2_2 [0]), .ZN(
        \Red_MCInst_MC2_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC2_v0_2 [0]), .B(\Red_MCInst_MC2_v1_2 [0]), .Z(\Red_MCInst_MC2_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC2_r2Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC2_r2Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[16]) );
  XNOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC2_v3_2 [1]), .B(\Red_MCInst_MC2_v2_2 [1]), .ZN(
        \Red_MCInst_MC2_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC2_v0_2 [1]), .B(\Red_MCInst_MC2_v1_2 [1]), .Z(\Red_MCInst_MC2_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC2_r2Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC2_r2Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[17]) );
  XNOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC2_v3_2 [2]), .B(\Red_MCInst_MC2_v2_2 [2]), .ZN(
        \Red_MCInst_MC2_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC2_v0_2 [2]), .B(\Red_MCInst_MC2_v1_2 [2]), .Z(\Red_MCInst_MC2_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC2_r3Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC2_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[3]) );
  XNOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC2_v3_3 [0]), .B(\Red_MCInst_MC2_v2_3 [0]), .ZN(
        \Red_MCInst_MC2_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC2_v0_3 [0]), .B(\Red_MCInst_MC2_v1_3 [0]), .Z(\Red_MCInst_MC2_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC2_r3Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC2_r3Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[4]) );
  XNOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC2_v3_3 [1]), .B(\Red_MCInst_MC2_v2_3 [1]), .ZN(
        \Red_MCInst_MC2_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC2_v0_3 [1]), .B(\Red_MCInst_MC2_v1_3 [1]), .Z(\Red_MCInst_MC2_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC2_r3Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC2_r3Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[5]) );
  XNOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC2_v3_3 [2]), .B(\Red_MCInst_MC2_v2_3 [2]), .ZN(
        \Red_MCInst_MC2_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC2_v0_3 [2]), .B(\Red_MCInst_MC2_v1_3 [2]), .Z(\Red_MCInst_MC2_r3Inst_XORInst_0_2_n5 ) );
  XOR2_X1 \Red_MCInst_MC3_v0_2Inst_0_U3  ( .A(\MCInst_MC3_v0_3 [3]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\Red_MCInst_MC3_v0_2 [0]) );
  XOR2_X1 \Red_MCInst_MC3_v0_3Inst_0_U3  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(
        \Red_MCInst_MC3_v0_2 [2]), .Z(\Red_MCInst_MC3_v0_3 [0]) );
  XNOR2_X1 \Red_MCInst_MC3_v1_0Inst_0_U4  ( .A(\Red_MCInst_MC3_v1_0Inst_0_n2 ), 
        .B(\Red_MCInst_MC3_v1_2 [1]), .ZN(\Red_MCInst_MC3_v1_0 [0]) );
  XNOR2_X1 \Red_MCInst_MC3_v1_0Inst_0_U3  ( .A(\MCInst_MC3_v1_3 [3]), .B(
        \MCInst_MC3_v1_0 [0]), .ZN(\Red_MCInst_MC3_v1_0Inst_0_n2 ) );
  XOR2_X1 \Red_MCInst_MC3_v1_2Inst_0_U3  ( .A(\Red_MCInst_MC3_v1_2 [1]), .B(
        \Red_MCInst_MC3_v1_1 [2]), .Z(\Red_MCInst_MC3_v1_2 [0]) );
  XOR2_X1 \Red_MCInst_MC3_v1_3Inst_0_U3  ( .A(\MCInst_MC3_v1_0 [0]), .B(
        \Red_MCInst_MC3_v1_2 [1]), .Z(\Red_MCInst_MC3_v1_3 [0]) );
  XOR2_X1 \Red_MCInst_MC3_v2_0Inst_0_U3  ( .A(\Red_MCInst_MC3_v2_1 [1]), .B(
        \MCInst_MC3_v2_0 [2]), .Z(\Red_MCInst_MC3_v2_0 [0]) );
  XOR2_X1 \Red_MCInst_MC3_v2_1Inst_0_U3  ( .A(\MCInst_MC3_v2_0 [2]), .B(
        \MCInst_MC3_v2_0 [3]), .Z(\Red_MCInst_MC3_v2_1 [0]) );
  XNOR2_X1 \Red_MCInst_MC3_v2_2Inst_0_U4  ( .A(\Red_MCInst_MC3_v2_2Inst_0_n2 ), 
        .B(\MCInst_MC3_v2_0 [2]), .ZN(\Red_MCInst_MC3_v2_2 [0]) );
  XNOR2_X1 \Red_MCInst_MC3_v2_2Inst_0_U3  ( .A(\Red_MCInst_MC3_v2_2 [1]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\Red_MCInst_MC3_v2_2Inst_0_n2 ) );
  XNOR2_X1 \Red_MCInst_MC3_v2_3Inst_0_U4  ( .A(\Red_MCInst_MC3_v2_3Inst_0_n2 ), 
        .B(\MCInst_MC3_v2_0 [3]), .ZN(\Red_MCInst_MC3_v2_3 [0]) );
  XNOR2_X1 \Red_MCInst_MC3_v2_3Inst_0_U3  ( .A(\Red_MCInst_MC3_v2_2 [1]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\Red_MCInst_MC3_v2_3Inst_0_n2 ) );
  XOR2_X1 \Red_MCInst_MC3_v3_0Inst_0_U3  ( .A(\MCInst_MC3_v3_2 [3]), .B(
        \Red_MCInst_MC3_v3_3 [2]), .Z(\Red_MCInst_MC3_v3_0 [0]) );
  XNOR2_X1 \Red_MCInst_MC3_v3_2Inst_0_U5  ( .A(\Red_MCInst_MC3_v3_2Inst_0_n4 ), 
        .B(\Red_MCInst_MC3_v3_2Inst_0_n3 ), .ZN(\Red_MCInst_MC3_v3_2 [0]) );
  XNOR2_X1 \Red_MCInst_MC3_v3_2Inst_0_U4  ( .A(\Red_MCInst_MC3_v3_3 [2]), .B(
        \MCInst_MC3_v3_2 [3]), .ZN(\Red_MCInst_MC3_v3_2Inst_0_n3 ) );
  XOR2_X1 \Red_MCInst_MC3_v3_2Inst_0_U3  ( .A(\MCInst_MC3_v3_0 [3]), .B(
        \Red_MCInst_MC3_v3_1 [2]), .Z(\Red_MCInst_MC3_v3_2Inst_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_v3_3Inst_0_U3  ( .A(\MCInst_MC3_v3_0 [3]), .B(
        \Red_MCInst_MC3_v3_1 [2]), .Z(\Red_MCInst_MC3_v3_3 [0]) );
  XOR2_X1 \Red_MCInst_MC3_v0_0Inst_1_U3  ( .A(\Red_MCInst_MC3_v0_2 [2]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\Red_MCInst_MC3_v0_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC3_v0_1Inst_1_U4  ( .A(\Red_MCInst_MC3_v0_1Inst_1_n2 ), 
        .B(\MCInst_MC3_v0_3 [3]), .ZN(\Red_MCInst_MC3_v0_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC3_v0_1Inst_1_U3  ( .A(\Red_MCInst_MC3_v0_1 [0]), .B(
        \Red_MCInst_MC3_v0_0 [0]), .ZN(\Red_MCInst_MC3_v0_1Inst_1_n2 ) );
  XOR2_X1 \Red_MCInst_MC3_v0_2Inst_1_U3  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(
        \Red_MCInst_MC3_v0_2 [2]), .Z(\Red_MCInst_MC3_v0_2 [1]) );
  XOR2_X1 \Red_MCInst_MC3_v0_3Inst_1_U3  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(
        \MCInst_MC3_v0_3 [3]), .Z(\Red_MCInst_MC3_v0_3 [1]) );
  XNOR2_X1 \Red_MCInst_MC3_v1_0Inst_1_U4  ( .A(\Red_MCInst_MC3_v1_0Inst_1_n2 ), 
        .B(\Red_MCInst_MC3_v1_2 [1]), .ZN(\Red_MCInst_MC3_v1_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC3_v1_0Inst_1_U3  ( .A(\Red_MCInst_MC3_v1_1 [2]), .B(
        \MCInst_MC3_v1_0 [0]), .ZN(\Red_MCInst_MC3_v1_0Inst_1_n2 ) );
  XNOR2_X1 \Red_MCInst_MC3_v1_1Inst_1_U5  ( .A(\Red_MCInst_MC3_v1_1Inst_1_n4 ), 
        .B(\Red_MCInst_MC3_v1_1Inst_1_n3 ), .ZN(\Red_MCInst_MC3_v1_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC3_v1_1Inst_1_U4  ( .A(\Red_MCInst_MC3_v1_2 [1]), .B(
        \MCInst_MC3_v1_0 [0]), .ZN(\Red_MCInst_MC3_v1_1Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_MC3_v1_1Inst_1_U3  ( .A(\MCInst_MC3_v1_3 [3]), .B(
        \Red_MCInst_MC3_v1_1 [2]), .Z(\Red_MCInst_MC3_v1_1Inst_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_v1_3Inst_1_U3  ( .A(\MCInst_MC3_v1_0 [0]), .B(
        \MCInst_MC3_v1_3 [3]), .Z(\Red_MCInst_MC3_v1_3 [1]) );
  XOR2_X1 \Red_MCInst_MC3_v2_0Inst_1_U3  ( .A(\Red_MCInst_MC3_v2_1 [1]), .B(
        \MCInst_MC3_v2_0 [3]), .Z(\Red_MCInst_MC3_v2_0 [1]) );
  XOR2_X1 \Red_MCInst_MC3_v2_3Inst_1_U3  ( .A(\Red_MCInst_MC3_v2_1 [1]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\Red_MCInst_MC3_v2_3 [1]) );
  XOR2_X1 \Red_MCInst_MC3_v3_0Inst_1_U3  ( .A(\MCInst_MC3_v3_2 [3]), .B(
        \MCInst_MC3_v3_0 [3]), .Z(\Red_MCInst_MC3_v3_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC3_v3_1Inst_1_U5  ( .A(\Red_MCInst_MC3_v3_1Inst_1_n4 ), 
        .B(\Red_MCInst_MC3_v3_1Inst_1_n3 ), .ZN(\Red_MCInst_MC3_v3_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC3_v3_1Inst_1_U4  ( .A(\Red_MCInst_MC3_v3_3 [2]), .B(
        \MCInst_MC3_v3_2 [3]), .ZN(\Red_MCInst_MC3_v3_1Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_MC3_v3_1Inst_1_U3  ( .A(\MCInst_MC3_v3_0 [3]), .B(
        \Red_MCInst_MC3_v3_1 [2]), .Z(\Red_MCInst_MC3_v3_1Inst_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_v3_2Inst_1_U3  ( .A(\Red_MCInst_MC3_v3_3 [2]), .B(
        \MCInst_MC3_v3_0 [3]), .Z(\Red_MCInst_MC3_v3_2 [1]) );
  XOR2_X1 \Red_MCInst_MC3_v3_3Inst_1_U3  ( .A(\MCInst_MC3_v3_2 [3]), .B(
        \Red_MCInst_MC3_v3_3 [2]), .Z(\Red_MCInst_MC3_v3_3 [1]) );
  XNOR2_X1 \Red_MCInst_MC3_v0_0Inst_2_U4  ( .A(\Red_MCInst_MC3_v0_0Inst_2_n2 ), 
        .B(\Red_MCInst_MC3_v0_2 [2]), .ZN(\Red_MCInst_MC3_v0_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v0_0Inst_2_U3  ( .A(\MCInst_MC3_v0_3 [3]), .B(
        \Red_MCInst_MC3_v0_0 [0]), .ZN(\Red_MCInst_MC3_v0_0Inst_2_n2 ) );
  XOR2_X1 \Red_MCInst_MC3_v0_1Inst_2_U3  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(
        \Red_MCInst_MC3_v0_2 [2]), .Z(\Red_MCInst_MC3_v0_1 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v0_3Inst_2_U5  ( .A(\Red_MCInst_MC3_v0_3Inst_2_n4 ), 
        .B(\Red_MCInst_MC3_v0_3Inst_2_n3 ), .ZN(\Red_MCInst_MC3_v0_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v0_3Inst_2_U4  ( .A(\Red_MCInst_MC3_v0_2 [2]), .B(
        \Red_MCInst_MC3_v0_0 [0]), .ZN(\Red_MCInst_MC3_v0_3Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC3_v0_3Inst_2_U3  ( .A(\MCInst_MC3_v0_3 [3]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\Red_MCInst_MC3_v0_3Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC3_v1_0Inst_2_U4  ( .A(\Red_MCInst_MC3_v1_0Inst_2_n2 ), 
        .B(\MCInst_MC3_v1_3 [3]), .ZN(\Red_MCInst_MC3_v1_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v1_0Inst_2_U3  ( .A(\Red_MCInst_MC3_v1_1 [2]), .B(
        \Red_MCInst_MC3_v1_2 [1]), .ZN(\Red_MCInst_MC3_v1_0Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC3_v1_2Inst_2_U4  ( .A(\Red_MCInst_MC3_v1_2Inst_2_n2 ), 
        .B(\Red_MCInst_MC3_v1_2 [1]), .ZN(\Red_MCInst_MC3_v1_2 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v1_2Inst_2_U3  ( .A(\Red_MCInst_MC3_v1_1 [2]), .B(
        \MCInst_MC3_v1_0 [0]), .ZN(\Red_MCInst_MC3_v1_2Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC3_v1_3Inst_2_U5  ( .A(\Red_MCInst_MC3_v1_3Inst_2_n4 ), 
        .B(\Red_MCInst_MC3_v1_3Inst_2_n3 ), .ZN(\Red_MCInst_MC3_v1_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v1_3Inst_2_U4  ( .A(\Red_MCInst_MC3_v1_2 [1]), .B(
        \MCInst_MC3_v1_0 [0]), .ZN(\Red_MCInst_MC3_v1_3Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC3_v1_3Inst_2_U3  ( .A(\MCInst_MC3_v1_3 [3]), .B(
        \Red_MCInst_MC3_v1_1 [2]), .Z(\Red_MCInst_MC3_v1_3Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC3_v2_0Inst_2_U5  ( .A(\Red_MCInst_MC3_v2_0Inst_2_n4 ), 
        .B(\Red_MCInst_MC3_v2_0Inst_2_n3 ), .ZN(\Red_MCInst_MC3_v2_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v2_0Inst_2_U4  ( .A(\MCInst_MC3_v2_0 [2]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\Red_MCInst_MC3_v2_0Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC3_v2_0Inst_2_U3  ( .A(\MCInst_MC3_v2_0 [3]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\Red_MCInst_MC3_v2_0Inst_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_v2_1Inst_2_U3  ( .A(\Red_MCInst_MC3_v2_1 [1]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\Red_MCInst_MC3_v2_1 [2]) );
  XOR2_X1 \Red_MCInst_MC3_v2_2Inst_2_U3  ( .A(\MCInst_MC3_v2_0 [3]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\Red_MCInst_MC3_v2_2 [2]) );
  XOR2_X1 \Red_MCInst_MC3_v2_3Inst_2_U3  ( .A(\Red_MCInst_MC3_v2_1 [1]), .B(
        \MCInst_MC3_v2_0 [3]), .Z(\Red_MCInst_MC3_v2_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v3_0Inst_2_U5  ( .A(\Red_MCInst_MC3_v3_0Inst_2_n4 ), 
        .B(\Red_MCInst_MC3_v3_0Inst_2_n3 ), .ZN(\Red_MCInst_MC3_v3_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v3_0Inst_2_U4  ( .A(\Red_MCInst_MC3_v3_3 [2]), .B(
        \MCInst_MC3_v3_2 [3]), .ZN(\Red_MCInst_MC3_v3_0Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC3_v3_0Inst_2_U3  ( .A(\MCInst_MC3_v3_0 [3]), .B(
        \Red_MCInst_MC3_v3_1 [2]), .Z(\Red_MCInst_MC3_v3_0Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC3_v3_2Inst_2_U4  ( .A(\Red_MCInst_MC3_v3_2Inst_2_n2 ), 
        .B(\MCInst_MC3_v3_0 [3]), .ZN(\Red_MCInst_MC3_v3_2 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v3_2Inst_2_U3  ( .A(\Red_MCInst_MC3_v3_1 [2]), .B(
        \MCInst_MC3_v3_2 [3]), .ZN(\Red_MCInst_MC3_v3_2Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC3_r0Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC3_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[36]) );
  XNOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC3_v3_0 [0]), .B(\Red_MCInst_MC3_v2_0 [0]), .ZN(
        \Red_MCInst_MC3_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(\Red_MCInst_MC3_v1_0 [0]), .Z(\Red_MCInst_MC3_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC3_r0Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC3_r0Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[37]) );
  XNOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC3_v3_0 [1]), .B(\Red_MCInst_MC3_v2_0 [1]), .ZN(
        \Red_MCInst_MC3_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC3_v0_0 [1]), .B(\Red_MCInst_MC3_v1_0 [1]), .Z(\Red_MCInst_MC3_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC3_r0Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC3_r0Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[38]) );
  XNOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC3_v3_0 [2]), .B(\Red_MCInst_MC3_v2_0 [2]), .ZN(
        \Red_MCInst_MC3_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC3_v0_0 [2]), .B(\Red_MCInst_MC3_v1_0 [2]), .Z(\Red_MCInst_MC3_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC3_r1Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC3_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[24]) );
  XNOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC3_v3_3 [2]), .B(\Red_MCInst_MC3_v2_1 [0]), .ZN(
        \Red_MCInst_MC3_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC3_v0_1 [0]), .B(\Red_MCInst_MC3_v1_2 [1]), .Z(\Red_MCInst_MC3_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC3_r1Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC3_r1Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[25]) );
  XNOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC3_v3_1 [1]), .B(\Red_MCInst_MC3_v2_1 [1]), .ZN(
        \Red_MCInst_MC3_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC3_v0_1 [1]), .B(\Red_MCInst_MC3_v1_1 [1]), .Z(\Red_MCInst_MC3_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC3_r1Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC3_r1Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[26]) );
  XNOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC3_v3_1 [2]), .B(\Red_MCInst_MC3_v2_1 [2]), .ZN(
        \Red_MCInst_MC3_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC3_v0_1 [2]), .B(\Red_MCInst_MC3_v1_1 [2]), .Z(\Red_MCInst_MC3_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC3_r2Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC3_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[12]) );
  XNOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC3_v3_2 [0]), .B(\Red_MCInst_MC3_v2_2 [0]), .ZN(
        \Red_MCInst_MC3_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC3_v0_2 [0]), .B(\Red_MCInst_MC3_v1_2 [0]), .Z(\Red_MCInst_MC3_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC3_r2Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC3_r2Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[13]) );
  XNOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC3_v3_2 [1]), .B(\Red_MCInst_MC3_v2_2 [1]), .ZN(
        \Red_MCInst_MC3_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC3_v0_2 [1]), .B(\Red_MCInst_MC3_v1_2 [1]), .Z(\Red_MCInst_MC3_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC3_r2Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC3_r2Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[14]) );
  XNOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC3_v3_2 [2]), .B(\Red_MCInst_MC3_v2_2 [2]), .ZN(
        \Red_MCInst_MC3_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC3_v0_2 [2]), .B(\Red_MCInst_MC3_v1_2 [2]), .Z(\Red_MCInst_MC3_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC3_r3Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC3_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[0]) );
  XNOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC3_v3_3 [0]), .B(\Red_MCInst_MC3_v2_3 [0]), .ZN(
        \Red_MCInst_MC3_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC3_v0_3 [0]), .B(\Red_MCInst_MC3_v1_3 [0]), .Z(\Red_MCInst_MC3_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC3_r3Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC3_r3Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[1]) );
  XNOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC3_v3_3 [1]), .B(\Red_MCInst_MC3_v2_3 [1]), .ZN(
        \Red_MCInst_MC3_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC3_v0_3 [1]), .B(\Red_MCInst_MC3_v1_3 [1]), .Z(\Red_MCInst_MC3_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC3_r3Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC3_r3Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[2]) );
  XNOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC3_v3_3 [2]), .B(\Red_MCInst_MC3_v2_3 [2]), .ZN(
        \Red_MCInst_MC3_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC3_v0_3 [2]), .B(\Red_MCInst_MC3_v1_3 [2]), .Z(\Red_MCInst_MC3_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_0_LFInst_0_n2 ), .B(StateRegOutput[1]), .ZN(
        Red_SignaltoCheck[0]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_0_U3  ( .A(StateRegOutput[2]), .B(
        StateRegOutput[0]), .ZN(\Red_ToCheckInst_LFInst_0_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_0_LFInst_1_n2 ), .B(StateRegOutput[1]), .ZN(
        Red_SignaltoCheck[1]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_1_U3  ( .A(StateRegOutput[3]), .B(
        StateRegOutput[0]), .ZN(\Red_ToCheckInst_LFInst_0_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_0_LFInst_2_n2 ), .B(StateRegOutput[2]), .ZN(
        Red_SignaltoCheck[2]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_2_U3  ( .A(StateRegOutput[3]), .B(
        StateRegOutput[1]), .ZN(\Red_ToCheckInst_LFInst_0_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_1_LFInst_0_n2 ), .B(StateRegOutput[5]), .ZN(
        Red_SignaltoCheck[3]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_0_U3  ( .A(StateRegOutput[6]), .B(
        StateRegOutput[4]), .ZN(\Red_ToCheckInst_LFInst_1_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_1_LFInst_1_n2 ), .B(StateRegOutput[5]), .ZN(
        Red_SignaltoCheck[4]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_1_U3  ( .A(StateRegOutput[7]), .B(
        StateRegOutput[4]), .ZN(\Red_ToCheckInst_LFInst_1_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_1_LFInst_2_n2 ), .B(StateRegOutput[6]), .ZN(
        Red_SignaltoCheck[5]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_2_U3  ( .A(StateRegOutput[7]), .B(
        StateRegOutput[5]), .ZN(\Red_ToCheckInst_LFInst_1_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_2_LFInst_0_n2 ), .B(AddConstOutput[1]), .ZN(
        Red_SignaltoCheck[6]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_0_U3  ( .A(AddConstOutput[2]), .B(
        AddConstOutput[0]), .ZN(\Red_ToCheckInst_LFInst_2_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_2_LFInst_1_n2 ), .B(AddConstOutput[1]), .ZN(
        Red_SignaltoCheck[7]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_1_U3  ( .A(AddConstOutput[3]), .B(
        AddConstOutput[0]), .ZN(\Red_ToCheckInst_LFInst_2_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_2_LFInst_2_n2 ), .B(AddConstOutput[2]), .ZN(
        Red_SignaltoCheck[8]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_2_U3  ( .A(AddConstOutput[3]), .B(
        AddConstOutput[1]), .ZN(\Red_ToCheckInst_LFInst_2_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_3_LFInst_0_n2 ), .B(AddConstOutput[5]), .ZN(
        Red_SignaltoCheck[9]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_0_U3  ( .A(AddConstOutput[6]), .B(
        AddConstOutput[4]), .ZN(\Red_ToCheckInst_LFInst_3_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_3_LFInst_1_n2 ), .B(AddConstOutput[5]), .ZN(
        Red_SignaltoCheck[10]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_1_U3  ( .A(AddConstOutput[7]), .B(
        AddConstOutput[4]), .ZN(\Red_ToCheckInst_LFInst_3_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_3_LFInst_2_n2 ), .B(AddConstOutput[6]), .ZN(
        Red_SignaltoCheck[11]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_2_U3  ( .A(AddConstOutput[7]), .B(
        AddConstOutput[5]), .ZN(\Red_ToCheckInst_LFInst_3_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_4_LFInst_0_n2 ), .B(StateRegOutput[17]), .ZN(
        Red_SignaltoCheck[12]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_0_U3  ( .A(StateRegOutput[18]), 
        .B(StateRegOutput[16]), .ZN(\Red_ToCheckInst_LFInst_4_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_4_LFInst_1_n2 ), .B(StateRegOutput[17]), .ZN(
        Red_SignaltoCheck[13]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_1_U3  ( .A(StateRegOutput[19]), 
        .B(StateRegOutput[16]), .ZN(\Red_ToCheckInst_LFInst_4_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_4_LFInst_2_n2 ), .B(StateRegOutput[18]), .ZN(
        Red_SignaltoCheck[14]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_2_U3  ( .A(StateRegOutput[19]), 
        .B(StateRegOutput[17]), .ZN(\Red_ToCheckInst_LFInst_4_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_5_LFInst_0_n2 ), .B(StateRegOutput[21]), .ZN(
        Red_SignaltoCheck[15]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_0_U3  ( .A(StateRegOutput[22]), 
        .B(StateRegOutput[20]), .ZN(\Red_ToCheckInst_LFInst_5_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_5_LFInst_1_n2 ), .B(StateRegOutput[21]), .ZN(
        Red_SignaltoCheck[16]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_1_U3  ( .A(StateRegOutput[23]), 
        .B(StateRegOutput[20]), .ZN(\Red_ToCheckInst_LFInst_5_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_5_LFInst_2_n2 ), .B(StateRegOutput[22]), .ZN(
        Red_SignaltoCheck[17]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_2_U3  ( .A(StateRegOutput[23]), 
        .B(StateRegOutput[21]), .ZN(\Red_ToCheckInst_LFInst_5_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_6_LFInst_0_n2 ), .B(AddConstOutput[9]), .ZN(
        Red_SignaltoCheck[18]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_0_U3  ( .A(AddConstOutput[10]), 
        .B(AddConstOutput[8]), .ZN(\Red_ToCheckInst_LFInst_6_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_6_LFInst_1_n2 ), .B(AddConstOutput[9]), .ZN(
        Red_SignaltoCheck[19]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_1_U3  ( .A(AddConstOutput[11]), 
        .B(AddConstOutput[8]), .ZN(\Red_ToCheckInst_LFInst_6_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_6_LFInst_2_n2 ), .B(AddConstOutput[10]), .ZN(
        Red_SignaltoCheck[20]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_2_U3  ( .A(AddConstOutput[11]), 
        .B(AddConstOutput[9]), .ZN(\Red_ToCheckInst_LFInst_6_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_7_LFInst_0_n2 ), .B(AddConstOutput[13]), .ZN(
        Red_SignaltoCheck[21]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_0_U3  ( .A(AddConstOutput[14]), 
        .B(AddConstOutput[12]), .ZN(\Red_ToCheckInst_LFInst_7_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_7_LFInst_1_n2 ), .B(AddConstOutput[13]), .ZN(
        Red_SignaltoCheck[22]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_1_U3  ( .A(AddConstOutput[15]), 
        .B(AddConstOutput[12]), .ZN(\Red_ToCheckInst_LFInst_7_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_7_LFInst_2_n2 ), .B(AddConstOutput[14]), .ZN(
        Red_SignaltoCheck[23]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_2_U3  ( .A(AddConstOutput[15]), 
        .B(AddConstOutput[13]), .ZN(\Red_ToCheckInst_LFInst_7_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_8_LFInst_0_n2 ), .B(StateRegOutput[33]), .ZN(
        Red_SignaltoCheck[24]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_0_U3  ( .A(StateRegOutput[34]), 
        .B(StateRegOutput[32]), .ZN(\Red_ToCheckInst_LFInst_8_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_8_LFInst_1_n2 ), .B(StateRegOutput[33]), .ZN(
        Red_SignaltoCheck[25]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_1_U3  ( .A(StateRegOutput[35]), 
        .B(StateRegOutput[32]), .ZN(\Red_ToCheckInst_LFInst_8_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_8_LFInst_2_n2 ), .B(StateRegOutput[34]), .ZN(
        Red_SignaltoCheck[26]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_2_U3  ( .A(StateRegOutput[35]), 
        .B(StateRegOutput[33]), .ZN(\Red_ToCheckInst_LFInst_8_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_9_LFInst_0_n2 ), .B(StateRegOutput[37]), .ZN(
        Red_SignaltoCheck[27]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_0_U3  ( .A(StateRegOutput[38]), 
        .B(StateRegOutput[36]), .ZN(\Red_ToCheckInst_LFInst_9_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_9_LFInst_1_n2 ), .B(StateRegOutput[37]), .ZN(
        Red_SignaltoCheck[28]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_1_U3  ( .A(StateRegOutput[39]), 
        .B(StateRegOutput[36]), .ZN(\Red_ToCheckInst_LFInst_9_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_9_LFInst_2_n2 ), .B(StateRegOutput[38]), .ZN(
        Red_SignaltoCheck[29]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_2_U3  ( .A(StateRegOutput[39]), 
        .B(StateRegOutput[37]), .ZN(\Red_ToCheckInst_LFInst_9_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_10_LFInst_0_n2 ), .B(AddConstOutput[17]), .ZN(
        Red_SignaltoCheck[30]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_0_U3  ( .A(AddConstOutput[18]), 
        .B(AddConstOutput[16]), .ZN(\Red_ToCheckInst_LFInst_10_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_10_LFInst_1_n2 ), .B(AddConstOutput[17]), .ZN(
        Red_SignaltoCheck[31]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_1_U3  ( .A(AddConstOutput[19]), 
        .B(AddConstOutput[16]), .ZN(\Red_ToCheckInst_LFInst_10_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_10_LFInst_2_n2 ), .B(AddConstOutput[18]), .ZN(
        Red_SignaltoCheck[32]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_2_U3  ( .A(AddConstOutput[19]), 
        .B(AddConstOutput[17]), .ZN(\Red_ToCheckInst_LFInst_10_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_11_LFInst_0_n2 ), .B(AddConstOutput[21]), .ZN(
        Red_SignaltoCheck[33]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_0_U3  ( .A(AddConstOutput[22]), 
        .B(AddConstOutput[20]), .ZN(\Red_ToCheckInst_LFInst_11_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_11_LFInst_1_n2 ), .B(AddConstOutput[21]), .ZN(
        Red_SignaltoCheck[34]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_1_U3  ( .A(AddConstOutput[23]), 
        .B(AddConstOutput[20]), .ZN(\Red_ToCheckInst_LFInst_11_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_11_LFInst_2_n2 ), .B(AddConstOutput[22]), .ZN(
        Red_SignaltoCheck[35]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_2_U3  ( .A(AddConstOutput[23]), 
        .B(AddConstOutput[21]), .ZN(\Red_ToCheckInst_LFInst_11_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_12_LFInst_0_n2 ), .B(StateRegOutput[49]), .ZN(
        Red_SignaltoCheck[36]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_0_U3  ( .A(StateRegOutput[50]), 
        .B(StateRegOutput[48]), .ZN(\Red_ToCheckInst_LFInst_12_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_12_LFInst_1_n2 ), .B(StateRegOutput[49]), .ZN(
        Red_SignaltoCheck[37]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_1_U3  ( .A(StateRegOutput[51]), 
        .B(StateRegOutput[48]), .ZN(\Red_ToCheckInst_LFInst_12_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_12_LFInst_2_n2 ), .B(StateRegOutput[50]), .ZN(
        Red_SignaltoCheck[38]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_2_U3  ( .A(StateRegOutput[51]), 
        .B(StateRegOutput[49]), .ZN(\Red_ToCheckInst_LFInst_12_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_13_LFInst_0_n2 ), .B(StateRegOutput[53]), .ZN(
        Red_SignaltoCheck[39]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_0_U3  ( .A(StateRegOutput[54]), 
        .B(StateRegOutput[52]), .ZN(\Red_ToCheckInst_LFInst_13_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_13_LFInst_1_n2 ), .B(StateRegOutput[53]), .ZN(
        Red_SignaltoCheck[40]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_1_U3  ( .A(StateRegOutput[55]), 
        .B(StateRegOutput[52]), .ZN(\Red_ToCheckInst_LFInst_13_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_13_LFInst_2_n2 ), .B(StateRegOutput[54]), .ZN(
        Red_SignaltoCheck[41]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_2_U3  ( .A(StateRegOutput[55]), 
        .B(StateRegOutput[53]), .ZN(\Red_ToCheckInst_LFInst_13_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_14_LFInst_0_n2 ), .B(AddConstOutput[25]), .ZN(
        Red_SignaltoCheck[42]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_0_U3  ( .A(AddConstOutput[26]), 
        .B(AddConstOutput[24]), .ZN(\Red_ToCheckInst_LFInst_14_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_14_LFInst_1_n2 ), .B(AddConstOutput[25]), .ZN(
        Red_SignaltoCheck[43]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_1_U3  ( .A(AddConstOutput[27]), 
        .B(AddConstOutput[24]), .ZN(\Red_ToCheckInst_LFInst_14_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_14_LFInst_2_n2 ), .B(AddConstOutput[26]), .ZN(
        Red_SignaltoCheck[44]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_2_U3  ( .A(AddConstOutput[27]), 
        .B(AddConstOutput[25]), .ZN(\Red_ToCheckInst_LFInst_14_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_15_LFInst_0_n2 ), .B(AddConstOutput[29]), .ZN(
        Red_SignaltoCheck[45]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_0_U3  ( .A(AddConstOutput[30]), 
        .B(AddConstOutput[28]), .ZN(\Red_ToCheckInst_LFInst_15_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_15_LFInst_1_n2 ), .B(AddConstOutput[29]), .ZN(
        Red_SignaltoCheck[46]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_1_U3  ( .A(AddConstOutput[31]), 
        .B(AddConstOutput[28]), .ZN(\Red_ToCheckInst_LFInst_15_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_15_LFInst_2_n2 ), .B(AddConstOutput[30]), .ZN(
        Red_SignaltoCheck[47]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_2_U3  ( .A(AddConstOutput[31]), 
        .B(AddConstOutput[29]), .ZN(\Red_ToCheckInst_LFInst_15_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_16_LFInst_0_n2 ), .B(Ciphertext[1]), .ZN(
        Red_SignaltoCheck[48]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_0_U3  ( .A(Ciphertext[2]), .B(
        Ciphertext[0]), .ZN(\Red_ToCheckInst_LFInst_16_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_16_LFInst_1_n2 ), .B(Ciphertext[1]), .ZN(
        Red_SignaltoCheck[49]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_1_U3  ( .A(Ciphertext[3]), .B(
        Ciphertext[0]), .ZN(\Red_ToCheckInst_LFInst_16_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_16_LFInst_2_n2 ), .B(Ciphertext[2]), .ZN(
        Red_SignaltoCheck[50]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_2_U3  ( .A(Ciphertext[3]), .B(
        Ciphertext[1]), .ZN(\Red_ToCheckInst_LFInst_16_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_17_LFInst_0_n2 ), .B(Ciphertext[5]), .ZN(
        Red_SignaltoCheck[51]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_0_U3  ( .A(Ciphertext[6]), .B(
        Ciphertext[4]), .ZN(\Red_ToCheckInst_LFInst_17_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_17_LFInst_1_n2 ), .B(Ciphertext[5]), .ZN(
        Red_SignaltoCheck[52]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_1_U3  ( .A(Ciphertext[7]), .B(
        Ciphertext[4]), .ZN(\Red_ToCheckInst_LFInst_17_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_17_LFInst_2_n2 ), .B(Ciphertext[6]), .ZN(
        Red_SignaltoCheck[53]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_2_U3  ( .A(Ciphertext[7]), .B(
        Ciphertext[5]), .ZN(\Red_ToCheckInst_LFInst_17_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_18_LFInst_0_n2 ), .B(Ciphertext[9]), .ZN(
        Red_SignaltoCheck[54]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_0_U3  ( .A(Ciphertext[10]), .B(
        Ciphertext[8]), .ZN(\Red_ToCheckInst_LFInst_18_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_18_LFInst_1_n2 ), .B(Ciphertext[9]), .ZN(
        Red_SignaltoCheck[55]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_1_U3  ( .A(Ciphertext[11]), .B(
        Ciphertext[8]), .ZN(\Red_ToCheckInst_LFInst_18_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_18_LFInst_2_n2 ), .B(Ciphertext[10]), .ZN(
        Red_SignaltoCheck[56]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_2_U3  ( .A(Ciphertext[11]), .B(
        Ciphertext[9]), .ZN(\Red_ToCheckInst_LFInst_18_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_19_LFInst_0_n2 ), .B(Ciphertext[13]), .ZN(
        Red_SignaltoCheck[57]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_0_U3  ( .A(Ciphertext[14]), .B(
        Ciphertext[12]), .ZN(\Red_ToCheckInst_LFInst_19_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_19_LFInst_1_n2 ), .B(Ciphertext[13]), .ZN(
        Red_SignaltoCheck[58]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_1_U3  ( .A(Ciphertext[15]), .B(
        Ciphertext[12]), .ZN(\Red_ToCheckInst_LFInst_19_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_19_LFInst_2_n2 ), .B(Ciphertext[14]), .ZN(
        Red_SignaltoCheck[59]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_2_U3  ( .A(Ciphertext[15]), .B(
        Ciphertext[13]), .ZN(\Red_ToCheckInst_LFInst_19_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_20_LFInst_0_n2 ), .B(Ciphertext[17]), .ZN(
        Red_SignaltoCheck[60]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_0_U3  ( .A(Ciphertext[18]), .B(
        Ciphertext[16]), .ZN(\Red_ToCheckInst_LFInst_20_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_20_LFInst_1_n2 ), .B(Ciphertext[17]), .ZN(
        Red_SignaltoCheck[61]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_1_U3  ( .A(Ciphertext[19]), .B(
        Ciphertext[16]), .ZN(\Red_ToCheckInst_LFInst_20_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_20_LFInst_2_n2 ), .B(Ciphertext[18]), .ZN(
        Red_SignaltoCheck[62]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_2_U3  ( .A(Ciphertext[19]), .B(
        Ciphertext[17]), .ZN(\Red_ToCheckInst_LFInst_20_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_21_LFInst_0_n2 ), .B(Ciphertext[21]), .ZN(
        Red_SignaltoCheck[63]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_0_U3  ( .A(Ciphertext[22]), .B(
        Ciphertext[20]), .ZN(\Red_ToCheckInst_LFInst_21_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_21_LFInst_1_n2 ), .B(Ciphertext[21]), .ZN(
        Red_SignaltoCheck[64]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_1_U3  ( .A(Ciphertext[23]), .B(
        Ciphertext[20]), .ZN(\Red_ToCheckInst_LFInst_21_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_21_LFInst_2_n2 ), .B(Ciphertext[22]), .ZN(
        Red_SignaltoCheck[65]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_2_U3  ( .A(Ciphertext[23]), .B(
        Ciphertext[21]), .ZN(\Red_ToCheckInst_LFInst_21_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_22_LFInst_0_n2 ), .B(Ciphertext[25]), .ZN(
        Red_SignaltoCheck[66]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_0_U3  ( .A(Ciphertext[26]), .B(
        Ciphertext[24]), .ZN(\Red_ToCheckInst_LFInst_22_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_22_LFInst_1_n2 ), .B(Ciphertext[25]), .ZN(
        Red_SignaltoCheck[67]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_1_U3  ( .A(Ciphertext[27]), .B(
        Ciphertext[24]), .ZN(\Red_ToCheckInst_LFInst_22_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_22_LFInst_2_n2 ), .B(Ciphertext[26]), .ZN(
        Red_SignaltoCheck[68]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_2_U3  ( .A(Ciphertext[27]), .B(
        Ciphertext[25]), .ZN(\Red_ToCheckInst_LFInst_22_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_23_LFInst_0_n2 ), .B(Ciphertext[29]), .ZN(
        Red_SignaltoCheck[69]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_0_U3  ( .A(Ciphertext[30]), .B(
        Ciphertext[28]), .ZN(\Red_ToCheckInst_LFInst_23_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_23_LFInst_1_n2 ), .B(Ciphertext[29]), .ZN(
        Red_SignaltoCheck[70]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_1_U3  ( .A(Ciphertext[31]), .B(
        Ciphertext[28]), .ZN(\Red_ToCheckInst_LFInst_23_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_23_LFInst_2_n2 ), .B(Ciphertext[30]), .ZN(
        Red_SignaltoCheck[71]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_2_U3  ( .A(Ciphertext[31]), .B(
        Ciphertext[29]), .ZN(\Red_ToCheckInst_LFInst_23_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_24_LFInst_0_n2 ), .B(Ciphertext[33]), .ZN(
        Red_SignaltoCheck[72]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_0_U3  ( .A(Ciphertext[34]), .B(
        Ciphertext[32]), .ZN(\Red_ToCheckInst_LFInst_24_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_24_LFInst_1_n2 ), .B(Ciphertext[33]), .ZN(
        Red_SignaltoCheck[73]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_1_U3  ( .A(Ciphertext[35]), .B(
        Ciphertext[32]), .ZN(\Red_ToCheckInst_LFInst_24_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_24_LFInst_2_n2 ), .B(Ciphertext[34]), .ZN(
        Red_SignaltoCheck[74]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_2_U3  ( .A(Ciphertext[35]), .B(
        Ciphertext[33]), .ZN(\Red_ToCheckInst_LFInst_24_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_25_LFInst_0_n2 ), .B(Ciphertext[37]), .ZN(
        Red_SignaltoCheck[75]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_0_U3  ( .A(Ciphertext[38]), .B(
        Ciphertext[36]), .ZN(\Red_ToCheckInst_LFInst_25_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_25_LFInst_1_n2 ), .B(Ciphertext[37]), .ZN(
        Red_SignaltoCheck[76]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_1_U3  ( .A(Ciphertext[39]), .B(
        Ciphertext[36]), .ZN(\Red_ToCheckInst_LFInst_25_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_25_LFInst_2_n2 ), .B(Ciphertext[38]), .ZN(
        Red_SignaltoCheck[77]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_2_U3  ( .A(Ciphertext[39]), .B(
        Ciphertext[37]), .ZN(\Red_ToCheckInst_LFInst_25_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_26_LFInst_0_n2 ), .B(Ciphertext[41]), .ZN(
        Red_SignaltoCheck[78]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_0_U3  ( .A(Ciphertext[42]), .B(
        Ciphertext[40]), .ZN(\Red_ToCheckInst_LFInst_26_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_26_LFInst_1_n2 ), .B(Ciphertext[41]), .ZN(
        Red_SignaltoCheck[79]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_1_U3  ( .A(Ciphertext[43]), .B(
        Ciphertext[40]), .ZN(\Red_ToCheckInst_LFInst_26_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_26_LFInst_2_n2 ), .B(Ciphertext[42]), .ZN(
        Red_SignaltoCheck[80]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_2_U3  ( .A(Ciphertext[43]), .B(
        Ciphertext[41]), .ZN(\Red_ToCheckInst_LFInst_26_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_27_LFInst_0_n2 ), .B(Ciphertext[45]), .ZN(
        Red_SignaltoCheck[81]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_0_U3  ( .A(Ciphertext[46]), .B(
        Ciphertext[44]), .ZN(\Red_ToCheckInst_LFInst_27_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_27_LFInst_1_n2 ), .B(Ciphertext[45]), .ZN(
        Red_SignaltoCheck[82]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_1_U3  ( .A(Ciphertext[47]), .B(
        Ciphertext[44]), .ZN(\Red_ToCheckInst_LFInst_27_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_27_LFInst_2_n2 ), .B(Ciphertext[46]), .ZN(
        Red_SignaltoCheck[83]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_2_U3  ( .A(Ciphertext[47]), .B(
        Ciphertext[45]), .ZN(\Red_ToCheckInst_LFInst_27_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_28_LFInst_0_n2 ), .B(Ciphertext[49]), .ZN(
        Red_SignaltoCheck[84]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_0_U3  ( .A(Ciphertext[50]), .B(
        Ciphertext[48]), .ZN(\Red_ToCheckInst_LFInst_28_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_28_LFInst_1_n2 ), .B(Ciphertext[49]), .ZN(
        Red_SignaltoCheck[85]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_1_U3  ( .A(Ciphertext[51]), .B(
        Ciphertext[48]), .ZN(\Red_ToCheckInst_LFInst_28_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_28_LFInst_2_n2 ), .B(Ciphertext[50]), .ZN(
        Red_SignaltoCheck[86]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_2_U3  ( .A(Ciphertext[51]), .B(
        Ciphertext[49]), .ZN(\Red_ToCheckInst_LFInst_28_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_29_LFInst_0_n2 ), .B(Ciphertext[53]), .ZN(
        Red_SignaltoCheck[87]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_0_U3  ( .A(Ciphertext[54]), .B(
        Ciphertext[52]), .ZN(\Red_ToCheckInst_LFInst_29_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_29_LFInst_1_n2 ), .B(Ciphertext[53]), .ZN(
        Red_SignaltoCheck[88]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_1_U3  ( .A(Ciphertext[55]), .B(
        Ciphertext[52]), .ZN(\Red_ToCheckInst_LFInst_29_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_29_LFInst_2_n2 ), .B(Ciphertext[54]), .ZN(
        Red_SignaltoCheck[89]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_2_U3  ( .A(Ciphertext[55]), .B(
        Ciphertext[53]), .ZN(\Red_ToCheckInst_LFInst_29_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_30_LFInst_0_n2 ), .B(Ciphertext[57]), .ZN(
        Red_SignaltoCheck[90]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_0_U3  ( .A(Ciphertext[58]), .B(
        Ciphertext[56]), .ZN(\Red_ToCheckInst_LFInst_30_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_30_LFInst_1_n2 ), .B(Ciphertext[57]), .ZN(
        Red_SignaltoCheck[91]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_1_U3  ( .A(Ciphertext[59]), .B(
        Ciphertext[56]), .ZN(\Red_ToCheckInst_LFInst_30_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_30_LFInst_2_n2 ), .B(Ciphertext[58]), .ZN(
        Red_SignaltoCheck[92]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_2_U3  ( .A(Ciphertext[59]), .B(
        Ciphertext[57]), .ZN(\Red_ToCheckInst_LFInst_30_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_31_LFInst_0_n2 ), .B(Ciphertext[61]), .ZN(
        Red_SignaltoCheck[93]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_0_U3  ( .A(Ciphertext[62]), .B(
        Ciphertext[60]), .ZN(\Red_ToCheckInst_LFInst_31_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_31_LFInst_1_n2 ), .B(Ciphertext[61]), .ZN(
        Red_SignaltoCheck[94]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_1_U3  ( .A(Ciphertext[63]), .B(
        Ciphertext[60]), .ZN(\Red_ToCheckInst_LFInst_31_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_31_LFInst_2_n2 ), .B(Ciphertext[62]), .ZN(
        Red_SignaltoCheck[95]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_2_U3  ( .A(Ciphertext[63]), .B(
        Ciphertext[61]), .ZN(\Red_ToCheckInst_LFInst_31_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_32_LFInst_0_n2 ), .B(\Red_MCInst_MC3_v3_3 [2]), 
        .ZN(Red_SignaltoCheck[96]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_0_U3  ( .A(\MCInst_MC3_v3_0 [3]), 
        .B(\MCInst_MC3_v3_2 [3]), .ZN(\Red_ToCheckInst_LFInst_32_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_32_LFInst_1_n2 ), .B(\Red_MCInst_MC3_v3_3 [2]), 
        .ZN(Red_SignaltoCheck[97]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_1_U3  ( .A(
        \Red_MCInst_MC3_v3_1 [2]), .B(\MCInst_MC3_v3_2 [3]), .ZN(
        \Red_ToCheckInst_LFInst_32_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_32_LFInst_2_n2 ), .B(\MCInst_MC3_v3_0 [3]), 
        .ZN(Red_SignaltoCheck[98]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_2_U3  ( .A(
        \Red_MCInst_MC3_v3_1 [2]), .B(\Red_MCInst_MC3_v3_3 [2]), .ZN(
        \Red_ToCheckInst_LFInst_32_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_33_LFInst_0_n2 ), .B(\Red_MCInst_MC2_v3_3 [2]), 
        .ZN(Red_SignaltoCheck[99]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_0_U3  ( .A(\MCInst_MC2_v3_0 [3]), 
        .B(\MCInst_MC2_v3_2 [3]), .ZN(\Red_ToCheckInst_LFInst_33_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_33_LFInst_1_n2 ), .B(\Red_MCInst_MC2_v3_3 [2]), 
        .ZN(Red_SignaltoCheck[100]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_1_U3  ( .A(
        \Red_MCInst_MC2_v3_1 [2]), .B(\MCInst_MC2_v3_2 [3]), .ZN(
        \Red_ToCheckInst_LFInst_33_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_33_LFInst_2_n2 ), .B(\MCInst_MC2_v3_0 [3]), 
        .ZN(Red_SignaltoCheck[101]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_2_U3  ( .A(
        \Red_MCInst_MC2_v3_1 [2]), .B(\Red_MCInst_MC2_v3_3 [2]), .ZN(
        \Red_ToCheckInst_LFInst_33_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_34_LFInst_0_n2 ), .B(\Red_MCInst_MC1_v3_3 [2]), 
        .ZN(Red_SignaltoCheck[102]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_0_U3  ( .A(\MCInst_MC1_v3_0 [3]), 
        .B(\MCInst_MC1_v3_2 [3]), .ZN(\Red_ToCheckInst_LFInst_34_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_34_LFInst_1_n2 ), .B(\Red_MCInst_MC1_v3_3 [2]), 
        .ZN(Red_SignaltoCheck[103]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_1_U3  ( .A(
        \Red_MCInst_MC1_v3_1 [2]), .B(\MCInst_MC1_v3_2 [3]), .ZN(
        \Red_ToCheckInst_LFInst_34_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_34_LFInst_2_n2 ), .B(\MCInst_MC1_v3_0 [3]), 
        .ZN(Red_SignaltoCheck[104]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_2_U3  ( .A(
        \Red_MCInst_MC1_v3_1 [2]), .B(\Red_MCInst_MC1_v3_3 [2]), .ZN(
        \Red_ToCheckInst_LFInst_34_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_35_LFInst_0_n2 ), .B(\Red_MCInst_MC0_v3_3 [2]), 
        .ZN(Red_SignaltoCheck[105]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_0_U3  ( .A(\MCInst_MC0_v3_0 [3]), 
        .B(\MCInst_MC0_v3_2 [3]), .ZN(\Red_ToCheckInst_LFInst_35_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_35_LFInst_1_n2 ), .B(\Red_MCInst_MC0_v3_3 [2]), 
        .ZN(Red_SignaltoCheck[106]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_1_U3  ( .A(
        \Red_MCInst_MC0_v3_1 [2]), .B(\MCInst_MC0_v3_2 [3]), .ZN(
        \Red_ToCheckInst_LFInst_35_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_35_LFInst_2_n2 ), .B(\MCInst_MC0_v3_0 [3]), 
        .ZN(Red_SignaltoCheck[107]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_2_U3  ( .A(
        \Red_MCInst_MC0_v3_1 [2]), .B(\Red_MCInst_MC0_v3_3 [2]), .ZN(
        \Red_ToCheckInst_LFInst_35_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_36_LFInst_0_n2 ), .B(\MCInst_MC3_v2_0 [2]), 
        .ZN(Red_SignaltoCheck[108]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_0_U3  ( .A(\MCInst_MC3_v2_0 [3]), 
        .B(\Red_MCInst_MC3_v2_1 [1]), .ZN(
        \Red_ToCheckInst_LFInst_36_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_36_LFInst_1_n2 ), .B(\MCInst_MC3_v2_0 [2]), 
        .ZN(Red_SignaltoCheck[109]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_1_U3  ( .A(
        \Red_MCInst_MC3_v2_2 [1]), .B(\Red_MCInst_MC3_v2_1 [1]), .ZN(
        \Red_ToCheckInst_LFInst_36_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_36_LFInst_2_n2 ), .B(\MCInst_MC3_v2_0 [3]), 
        .ZN(Red_SignaltoCheck[110]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_2_U3  ( .A(
        \Red_MCInst_MC3_v2_2 [1]), .B(\MCInst_MC3_v2_0 [2]), .ZN(
        \Red_ToCheckInst_LFInst_36_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_37_LFInst_0_n2 ), .B(\MCInst_MC2_v2_0 [2]), 
        .ZN(Red_SignaltoCheck[111]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_0_U3  ( .A(\MCInst_MC2_v2_0 [3]), 
        .B(\Red_MCInst_MC2_v2_1 [1]), .ZN(
        \Red_ToCheckInst_LFInst_37_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_37_LFInst_1_n2 ), .B(\MCInst_MC2_v2_0 [2]), 
        .ZN(Red_SignaltoCheck[112]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_1_U3  ( .A(
        \Red_MCInst_MC2_v2_2 [1]), .B(\Red_MCInst_MC2_v2_1 [1]), .ZN(
        \Red_ToCheckInst_LFInst_37_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_37_LFInst_2_n2 ), .B(\MCInst_MC2_v2_0 [3]), 
        .ZN(Red_SignaltoCheck[113]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_2_U3  ( .A(
        \Red_MCInst_MC2_v2_2 [1]), .B(\MCInst_MC2_v2_0 [2]), .ZN(
        \Red_ToCheckInst_LFInst_37_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_38_LFInst_0_n2 ), .B(\MCInst_MC1_v2_0 [2]), 
        .ZN(Red_SignaltoCheck[114]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_0_U3  ( .A(\MCInst_MC1_v2_0 [3]), 
        .B(\Red_MCInst_MC1_v2_1 [1]), .ZN(
        \Red_ToCheckInst_LFInst_38_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_38_LFInst_1_n2 ), .B(\MCInst_MC1_v2_0 [2]), 
        .ZN(Red_SignaltoCheck[115]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_1_U3  ( .A(
        \Red_MCInst_MC1_v2_2 [1]), .B(\Red_MCInst_MC1_v2_1 [1]), .ZN(
        \Red_ToCheckInst_LFInst_38_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_38_LFInst_2_n2 ), .B(\MCInst_MC1_v2_0 [3]), 
        .ZN(Red_SignaltoCheck[116]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_2_U3  ( .A(
        \Red_MCInst_MC1_v2_2 [1]), .B(\MCInst_MC1_v2_0 [2]), .ZN(
        \Red_ToCheckInst_LFInst_38_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_39_LFInst_0_n2 ), .B(\MCInst_MC0_v2_0 [2]), 
        .ZN(Red_SignaltoCheck[117]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_0_U3  ( .A(\MCInst_MC0_v2_0 [3]), 
        .B(\Red_MCInst_MC0_v2_1 [1]), .ZN(
        \Red_ToCheckInst_LFInst_39_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_39_LFInst_1_n2 ), .B(\MCInst_MC0_v2_0 [2]), 
        .ZN(Red_SignaltoCheck[118]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_1_U3  ( .A(
        \Red_MCInst_MC0_v2_2 [1]), .B(\Red_MCInst_MC0_v2_1 [1]), .ZN(
        \Red_ToCheckInst_LFInst_39_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_39_LFInst_2_n2 ), .B(\MCInst_MC0_v2_0 [3]), 
        .ZN(Red_SignaltoCheck[119]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_2_U3  ( .A(
        \Red_MCInst_MC0_v2_2 [1]), .B(\MCInst_MC0_v2_0 [2]), .ZN(
        \Red_ToCheckInst_LFInst_39_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_40_LFInst_0_n2 ), .B(\Red_MCInst_MC3_v1_2 [1]), 
        .ZN(Red_SignaltoCheck[120]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_0_U3  ( .A(\MCInst_MC3_v1_3 [3]), 
        .B(\MCInst_MC3_v1_0 [0]), .ZN(\Red_ToCheckInst_LFInst_40_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_40_LFInst_1_n2 ), .B(\Red_MCInst_MC3_v1_2 [1]), 
        .ZN(Red_SignaltoCheck[121]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_1_U3  ( .A(
        \Red_MCInst_MC3_v1_1 [2]), .B(\MCInst_MC3_v1_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_40_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_40_LFInst_2_n2 ), .B(\MCInst_MC3_v1_3 [3]), 
        .ZN(Red_SignaltoCheck[122]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_2_U3  ( .A(
        \Red_MCInst_MC3_v1_1 [2]), .B(\Red_MCInst_MC3_v1_2 [1]), .ZN(
        \Red_ToCheckInst_LFInst_40_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_41_LFInst_0_n2 ), .B(\Red_MCInst_MC2_v1_2 [1]), 
        .ZN(Red_SignaltoCheck[123]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_0_U3  ( .A(\MCInst_MC2_v1_3 [3]), 
        .B(\MCInst_MC2_v1_0 [0]), .ZN(\Red_ToCheckInst_LFInst_41_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_41_LFInst_1_n2 ), .B(\Red_MCInst_MC2_v1_2 [1]), 
        .ZN(Red_SignaltoCheck[124]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_1_U3  ( .A(
        \Red_MCInst_MC2_v1_1 [2]), .B(\MCInst_MC2_v1_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_41_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_41_LFInst_2_n2 ), .B(\MCInst_MC2_v1_3 [3]), 
        .ZN(Red_SignaltoCheck[125]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_2_U3  ( .A(
        \Red_MCInst_MC2_v1_1 [2]), .B(\Red_MCInst_MC2_v1_2 [1]), .ZN(
        \Red_ToCheckInst_LFInst_41_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_42_LFInst_0_n2 ), .B(\Red_MCInst_MC1_v1_2 [1]), 
        .ZN(Red_SignaltoCheck[126]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_0_U3  ( .A(\MCInst_MC1_v1_3 [3]), 
        .B(\MCInst_MC1_v1_0 [0]), .ZN(\Red_ToCheckInst_LFInst_42_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_42_LFInst_1_n2 ), .B(\Red_MCInst_MC1_v1_2 [1]), 
        .ZN(Red_SignaltoCheck[127]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_1_U3  ( .A(
        \Red_MCInst_MC1_v1_1 [2]), .B(\MCInst_MC1_v1_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_42_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_42_LFInst_2_n2 ), .B(\MCInst_MC1_v1_3 [3]), 
        .ZN(Red_SignaltoCheck[128]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_2_U3  ( .A(
        \Red_MCInst_MC1_v1_1 [2]), .B(\Red_MCInst_MC1_v1_2 [1]), .ZN(
        \Red_ToCheckInst_LFInst_42_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_43_LFInst_0_n2 ), .B(\Red_MCInst_MC0_v1_2 [1]), 
        .ZN(Red_SignaltoCheck[129]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_0_U3  ( .A(\MCInst_MC0_v1_3 [3]), 
        .B(\MCInst_MC0_v1_0 [0]), .ZN(\Red_ToCheckInst_LFInst_43_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_43_LFInst_1_n2 ), .B(\Red_MCInst_MC0_v1_2 [1]), 
        .ZN(Red_SignaltoCheck[130]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_1_U3  ( .A(
        \Red_MCInst_MC0_v1_1 [2]), .B(\MCInst_MC0_v1_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_43_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_43_LFInst_2_n2 ), .B(\MCInst_MC0_v1_3 [3]), 
        .ZN(Red_SignaltoCheck[131]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_2_U3  ( .A(
        \Red_MCInst_MC0_v1_1 [2]), .B(\Red_MCInst_MC0_v1_2 [1]), .ZN(
        \Red_ToCheckInst_LFInst_43_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_44_LFInst_0_n2 ), .B(\Red_MCInst_MC3_v0_2 [2]), 
        .ZN(Red_SignaltoCheck[132]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_0_U3  ( .A(\MCInst_MC3_v0_3 [3]), 
        .B(\Red_MCInst_MC3_v0_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_44_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_44_LFInst_1_n2 ), .B(\Red_MCInst_MC3_v0_2 [2]), 
        .ZN(Red_SignaltoCheck[133]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_1_U3  ( .A(
        \Red_MCInst_MC3_v0_1 [0]), .B(\Red_MCInst_MC3_v0_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_44_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_44_LFInst_2_n2 ), .B(\MCInst_MC3_v0_3 [3]), 
        .ZN(Red_SignaltoCheck[134]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_2_U3  ( .A(
        \Red_MCInst_MC3_v0_1 [0]), .B(\Red_MCInst_MC3_v0_2 [2]), .ZN(
        \Red_ToCheckInst_LFInst_44_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_45_LFInst_0_n2 ), .B(\Red_MCInst_MC2_v0_2 [2]), 
        .ZN(Red_SignaltoCheck[135]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_0_U3  ( .A(\MCInst_MC2_v0_3 [3]), 
        .B(\Red_MCInst_MC2_v0_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_45_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_45_LFInst_1_n2 ), .B(\Red_MCInst_MC2_v0_2 [2]), 
        .ZN(Red_SignaltoCheck[136]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_1_U3  ( .A(
        \Red_MCInst_MC2_v0_1 [0]), .B(\Red_MCInst_MC2_v0_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_45_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_45_LFInst_2_n2 ), .B(\MCInst_MC2_v0_3 [3]), 
        .ZN(Red_SignaltoCheck[137]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_2_U3  ( .A(
        \Red_MCInst_MC2_v0_1 [0]), .B(\Red_MCInst_MC2_v0_2 [2]), .ZN(
        \Red_ToCheckInst_LFInst_45_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_46_LFInst_0_n2 ), .B(\Red_MCInst_MC1_v0_2 [2]), 
        .ZN(Red_SignaltoCheck[138]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_0_U3  ( .A(\MCInst_MC1_v0_3 [3]), 
        .B(\Red_MCInst_MC1_v0_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_46_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_46_LFInst_1_n2 ), .B(\Red_MCInst_MC1_v0_2 [2]), 
        .ZN(Red_SignaltoCheck[139]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_1_U3  ( .A(
        \Red_MCInst_MC1_v0_1 [0]), .B(\Red_MCInst_MC1_v0_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_46_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_46_LFInst_2_n2 ), .B(\MCInst_MC1_v0_3 [3]), 
        .ZN(Red_SignaltoCheck[140]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_2_U3  ( .A(
        \Red_MCInst_MC1_v0_1 [0]), .B(\Red_MCInst_MC1_v0_2 [2]), .ZN(
        \Red_ToCheckInst_LFInst_46_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_47_LFInst_0_n2 ), .B(\Red_MCInst_MC0_v0_2 [2]), 
        .ZN(Red_SignaltoCheck[141]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_0_U3  ( .A(\MCInst_MC0_v0_3 [3]), 
        .B(\Red_MCInst_MC0_v0_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_47_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_47_LFInst_1_n2 ), .B(\Red_MCInst_MC0_v0_2 [2]), 
        .ZN(Red_SignaltoCheck[142]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_1_U3  ( .A(
        \Red_MCInst_MC0_v0_1 [0]), .B(\Red_MCInst_MC0_v0_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_47_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_47_LFInst_2_n2 ), .B(\MCInst_MC0_v0_3 [3]), 
        .ZN(Red_SignaltoCheck[143]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_2_U3  ( .A(
        \Red_MCInst_MC0_v0_1 [0]), .B(\Red_MCInst_MC0_v0_2 [2]), .ZN(
        \Red_ToCheckInst_LFInst_47_LFInst_2_n2 ) );
  NOR2_X1 \Check1_CheckInst_0_U95  ( .A1(\Check1_CheckInst_0_n94 ), .A2(
        \Check1_CheckInst_0_n93 ), .ZN(Error[0]) );
  NAND2_X1 \Check1_CheckInst_0_U94  ( .A1(\Check1_CheckInst_0_n92 ), .A2(
        \Check1_CheckInst_0_n91 ), .ZN(\Check1_CheckInst_0_n93 ) );
  NOR2_X1 \Check1_CheckInst_0_U93  ( .A1(\Check1_CheckInst_0_n90 ), .A2(
        \Check1_CheckInst_0_n89 ), .ZN(\Check1_CheckInst_0_n91 ) );
  NAND2_X1 \Check1_CheckInst_0_U92  ( .A1(\Check1_CheckInst_0_n88 ), .A2(
        \Check1_CheckInst_0_n87 ), .ZN(\Check1_CheckInst_0_n89 ) );
  NOR2_X1 \Check1_CheckInst_0_U91  ( .A1(\Check1_CheckInst_0_n86 ), .A2(
        \Check1_CheckInst_0_n85 ), .ZN(\Check1_CheckInst_0_n87 ) );
  NAND2_X1 \Check1_CheckInst_0_U90  ( .A1(\Check1_CheckInst_0_n84 ), .A2(
        \Check1_CheckInst_0_n83 ), .ZN(\Check1_CheckInst_0_n85 ) );
  NOR2_X1 \Check1_CheckInst_0_U89  ( .A1(\Check1_CheckInst_0_n82 ), .A2(
        \Check1_CheckInst_0_n81 ), .ZN(\Check1_CheckInst_0_n83 ) );
  NAND2_X1 \Check1_CheckInst_0_U88  ( .A1(\Check1_CheckInst_0_n80 ), .A2(
        \Check1_CheckInst_0_n79 ), .ZN(\Check1_CheckInst_0_n81 ) );
  XNOR2_X1 \Check1_CheckInst_0_U87  ( .A(Red_ShiftRowsOutput[18]), .B(
        Red_SignaltoCheck[114]), .ZN(\Check1_CheckInst_0_n79 ) );
  XNOR2_X1 \Check1_CheckInst_0_U86  ( .A(Red_ShiftRowsOutput[21]), .B(
        Red_SignaltoCheck[117]), .ZN(\Check1_CheckInst_0_n80 ) );
  NAND2_X1 \Check1_CheckInst_0_U85  ( .A1(\Check1_CheckInst_0_n78 ), .A2(
        \Check1_CheckInst_0_n77 ), .ZN(\Check1_CheckInst_0_n82 ) );
  XNOR2_X1 \Check1_CheckInst_0_U84  ( .A(Red_ShiftRowsOutput[33]), .B(
        Red_SignaltoCheck[129]), .ZN(\Check1_CheckInst_0_n77 ) );
  XNOR2_X1 \Check1_CheckInst_0_U83  ( .A(Red_ShiftRowsOutput[27]), .B(
        Red_SignaltoCheck[123]), .ZN(\Check1_CheckInst_0_n78 ) );
  NOR2_X1 \Check1_CheckInst_0_U82  ( .A1(\Check1_CheckInst_0_n76 ), .A2(
        \Check1_CheckInst_0_n75 ), .ZN(\Check1_CheckInst_0_n84 ) );
  NAND2_X1 \Check1_CheckInst_0_U81  ( .A1(\Check1_CheckInst_0_n74 ), .A2(
        \Check1_CheckInst_0_n73 ), .ZN(\Check1_CheckInst_0_n75 ) );
  XNOR2_X1 \Check1_CheckInst_0_U80  ( .A(Red_ShiftRowsOutput[15]), .B(
        Red_SignaltoCheck[111]), .ZN(\Check1_CheckInst_0_n73 ) );
  XNOR2_X1 \Check1_CheckInst_0_U79  ( .A(Red_ShiftRowsOutput[9]), .B(
        Red_SignaltoCheck[105]), .ZN(\Check1_CheckInst_0_n74 ) );
  NAND2_X1 \Check1_CheckInst_0_U78  ( .A1(\Check1_CheckInst_0_n72 ), .A2(
        \Check1_CheckInst_0_n71 ), .ZN(\Check1_CheckInst_0_n76 ) );
  XNOR2_X1 \Check1_CheckInst_0_U77  ( .A(Red_ShiftRowsOutput[12]), .B(
        Red_SignaltoCheck[108]), .ZN(\Check1_CheckInst_0_n71 ) );
  XNOR2_X1 \Check1_CheckInst_0_U76  ( .A(Red_ShiftRowsOutput[24]), .B(
        Red_SignaltoCheck[120]), .ZN(\Check1_CheckInst_0_n72 ) );
  NAND2_X1 \Check1_CheckInst_0_U75  ( .A1(\Check1_CheckInst_0_n70 ), .A2(
        \Check1_CheckInst_0_n69 ), .ZN(\Check1_CheckInst_0_n86 ) );
  NOR2_X1 \Check1_CheckInst_0_U74  ( .A1(\Check1_CheckInst_0_n68 ), .A2(
        \Check1_CheckInst_0_n67 ), .ZN(\Check1_CheckInst_0_n69 ) );
  XOR2_X1 \Check1_CheckInst_0_U73  ( .A(Red_AddConstOutput[6]), .B(
        Red_SignaltoCheck[18]), .Z(\Check1_CheckInst_0_n67 ) );
  XOR2_X1 \Check1_CheckInst_0_U72  ( .A(Red_AddConstOutput[12]), .B(
        Red_SignaltoCheck[30]), .Z(\Check1_CheckInst_0_n68 ) );
  NOR2_X1 \Check1_CheckInst_0_U71  ( .A1(\Check1_CheckInst_0_n66 ), .A2(
        \Check1_CheckInst_0_n65 ), .ZN(\Check1_CheckInst_0_n70 ) );
  XOR2_X1 \Check1_CheckInst_0_U70  ( .A(Red_StateRegOutput[24]), .B(
        Red_SignaltoCheck[24]), .Z(\Check1_CheckInst_0_n65 ) );
  XOR2_X1 \Check1_CheckInst_0_U69  ( .A(Red_StateRegOutput[27]), .B(
        Red_SignaltoCheck[27]), .Z(\Check1_CheckInst_0_n66 ) );
  NOR2_X1 \Check1_CheckInst_0_U68  ( .A1(\Check1_CheckInst_0_n64 ), .A2(
        \Check1_CheckInst_0_n63 ), .ZN(\Check1_CheckInst_0_n88 ) );
  NAND2_X1 \Check1_CheckInst_0_U67  ( .A1(\Check1_CheckInst_0_n62 ), .A2(
        \Check1_CheckInst_0_n61 ), .ZN(\Check1_CheckInst_0_n63 ) );
  XNOR2_X1 \Check1_CheckInst_0_U66  ( .A(Red_AddConstOutput[0]), .B(
        Red_SignaltoCheck[6]), .ZN(\Check1_CheckInst_0_n61 ) );
  XNOR2_X1 \Check1_CheckInst_0_U65  ( .A(Red_AddConstOutput[3]), .B(
        Red_SignaltoCheck[9]), .ZN(\Check1_CheckInst_0_n62 ) );
  NAND2_X1 \Check1_CheckInst_0_U64  ( .A1(\Check1_CheckInst_0_n60 ), .A2(
        \Check1_CheckInst_0_n59 ), .ZN(\Check1_CheckInst_0_n64 ) );
  XNOR2_X1 \Check1_CheckInst_0_U63  ( .A(Red_AddConstOutput[9]), .B(
        Red_SignaltoCheck[21]), .ZN(\Check1_CheckInst_0_n59 ) );
  XNOR2_X1 \Check1_CheckInst_0_U62  ( .A(Red_StateRegOutput[15]), .B(
        Red_SignaltoCheck[15]), .ZN(\Check1_CheckInst_0_n60 ) );
  NAND2_X1 \Check1_CheckInst_0_U61  ( .A1(\Check1_CheckInst_0_n58 ), .A2(
        \Check1_CheckInst_0_n57 ), .ZN(\Check1_CheckInst_0_n90 ) );
  NOR2_X1 \Check1_CheckInst_0_U60  ( .A1(\Check1_CheckInst_0_n56 ), .A2(
        \Check1_CheckInst_0_n55 ), .ZN(\Check1_CheckInst_0_n57 ) );
  NAND2_X1 \Check1_CheckInst_0_U59  ( .A1(\Check1_CheckInst_0_n54 ), .A2(
        \Check1_CheckInst_0_n53 ), .ZN(\Check1_CheckInst_0_n55 ) );
  NOR2_X1 \Check1_CheckInst_0_U58  ( .A1(\Check1_CheckInst_0_n52 ), .A2(
        \Check1_CheckInst_0_n51 ), .ZN(\Check1_CheckInst_0_n53 ) );
  NAND2_X1 \Check1_CheckInst_0_U57  ( .A1(\Check1_CheckInst_0_n50 ), .A2(
        \Check1_CheckInst_0_n49 ), .ZN(\Check1_CheckInst_0_n51 ) );
  XNOR2_X1 \Check1_CheckInst_0_U56  ( .A(Red_ShiftRowsOutput[45]), .B(
        Red_SignaltoCheck[141]), .ZN(\Check1_CheckInst_0_n49 ) );
  XNOR2_X1 \Check1_CheckInst_0_U55  ( .A(Red_SignaltoCheck[3]), .B(
        Red_StateRegOutput[3]), .ZN(\Check1_CheckInst_0_n50 ) );
  NAND2_X1 \Check1_CheckInst_0_U54  ( .A1(\Check1_CheckInst_0_n48 ), .A2(
        \Check1_CheckInst_0_n47 ), .ZN(\Check1_CheckInst_0_n52 ) );
  XNOR2_X1 \Check1_CheckInst_0_U53  ( .A(Red_StateRegOutput[0]), .B(
        Red_SignaltoCheck[0]), .ZN(\Check1_CheckInst_0_n47 ) );
  XNOR2_X1 \Check1_CheckInst_0_U52  ( .A(Red_StateRegOutput[12]), .B(
        Red_SignaltoCheck[12]), .ZN(\Check1_CheckInst_0_n48 ) );
  NOR2_X1 \Check1_CheckInst_0_U51  ( .A1(\Check1_CheckInst_0_n46 ), .A2(
        \Check1_CheckInst_0_n45 ), .ZN(\Check1_CheckInst_0_n54 ) );
  NAND2_X1 \Check1_CheckInst_0_U50  ( .A1(\Check1_CheckInst_0_n44 ), .A2(
        \Check1_CheckInst_0_n43 ), .ZN(\Check1_CheckInst_0_n45 ) );
  XNOR2_X1 \Check1_CheckInst_0_U49  ( .A(Red_Feedback[6]), .B(
        Red_SignaltoCheck[54]), .ZN(\Check1_CheckInst_0_n43 ) );
  XNOR2_X1 \Check1_CheckInst_0_U48  ( .A(Red_Feedback[18]), .B(
        Red_SignaltoCheck[66]), .ZN(\Check1_CheckInst_0_n44 ) );
  NAND2_X1 \Check1_CheckInst_0_U47  ( .A1(\Check1_CheckInst_0_n42 ), .A2(
        \Check1_CheckInst_0_n41 ), .ZN(\Check1_CheckInst_0_n46 ) );
  XNOR2_X1 \Check1_CheckInst_0_U46  ( .A(Red_Feedback[12]), .B(
        Red_SignaltoCheck[60]), .ZN(\Check1_CheckInst_0_n41 ) );
  XNOR2_X1 \Check1_CheckInst_0_U45  ( .A(Red_Feedback[15]), .B(
        Red_SignaltoCheck[63]), .ZN(\Check1_CheckInst_0_n42 ) );
  NAND2_X1 \Check1_CheckInst_0_U44  ( .A1(\Check1_CheckInst_0_n40 ), .A2(
        \Check1_CheckInst_0_n39 ), .ZN(\Check1_CheckInst_0_n56 ) );
  NOR2_X1 \Check1_CheckInst_0_U43  ( .A1(\Check1_CheckInst_0_n38 ), .A2(
        \Check1_CheckInst_0_n37 ), .ZN(\Check1_CheckInst_0_n39 ) );
  XOR2_X1 \Check1_CheckInst_0_U42  ( .A(Red_AddConstOutput[18]), .B(
        Red_SignaltoCheck[42]), .Z(\Check1_CheckInst_0_n37 ) );
  XOR2_X1 \Check1_CheckInst_0_U41  ( .A(Red_AddConstOutput[21]), .B(
        Red_SignaltoCheck[45]), .Z(\Check1_CheckInst_0_n38 ) );
  NOR2_X1 \Check1_CheckInst_0_U40  ( .A1(\Check1_CheckInst_0_n36 ), .A2(
        \Check1_CheckInst_0_n35 ), .ZN(\Check1_CheckInst_0_n40 ) );
  XOR2_X1 \Check1_CheckInst_0_U39  ( .A(Red_Feedback[9]), .B(
        Red_SignaltoCheck[57]), .Z(\Check1_CheckInst_0_n35 ) );
  XOR2_X1 \Check1_CheckInst_0_U38  ( .A(Red_Feedback[3]), .B(
        Red_SignaltoCheck[51]), .Z(\Check1_CheckInst_0_n36 ) );
  NOR2_X1 \Check1_CheckInst_0_U37  ( .A1(\Check1_CheckInst_0_n34 ), .A2(
        \Check1_CheckInst_0_n33 ), .ZN(\Check1_CheckInst_0_n58 ) );
  NAND2_X1 \Check1_CheckInst_0_U36  ( .A1(\Check1_CheckInst_0_n32 ), .A2(
        \Check1_CheckInst_0_n31 ), .ZN(\Check1_CheckInst_0_n33 ) );
  XNOR2_X1 \Check1_CheckInst_0_U35  ( .A(Red_StateRegOutput[39]), .B(
        Red_SignaltoCheck[39]), .ZN(\Check1_CheckInst_0_n31 ) );
  XNOR2_X1 \Check1_CheckInst_0_U34  ( .A(Red_AddConstOutput[15]), .B(
        Red_SignaltoCheck[33]), .ZN(\Check1_CheckInst_0_n32 ) );
  NAND2_X1 \Check1_CheckInst_0_U33  ( .A1(\Check1_CheckInst_0_n30 ), .A2(
        \Check1_CheckInst_0_n29 ), .ZN(\Check1_CheckInst_0_n34 ) );
  XNOR2_X1 \Check1_CheckInst_0_U32  ( .A(Red_StateRegOutput[36]), .B(
        Red_SignaltoCheck[36]), .ZN(\Check1_CheckInst_0_n29 ) );
  XNOR2_X1 \Check1_CheckInst_0_U31  ( .A(Red_Feedback[0]), .B(
        Red_SignaltoCheck[48]), .ZN(\Check1_CheckInst_0_n30 ) );
  NOR2_X1 \Check1_CheckInst_0_U30  ( .A1(\Check1_CheckInst_0_n28 ), .A2(
        \Check1_CheckInst_0_n27 ), .ZN(\Check1_CheckInst_0_n92 ) );
  NAND2_X1 \Check1_CheckInst_0_U29  ( .A1(\Check1_CheckInst_0_n26 ), .A2(
        \Check1_CheckInst_0_n25 ), .ZN(\Check1_CheckInst_0_n27 ) );
  NOR2_X1 \Check1_CheckInst_0_U28  ( .A1(\Check1_CheckInst_0_n24 ), .A2(
        \Check1_CheckInst_0_n23 ), .ZN(\Check1_CheckInst_0_n25 ) );
  NAND2_X1 \Check1_CheckInst_0_U27  ( .A1(\Check1_CheckInst_0_n22 ), .A2(
        \Check1_CheckInst_0_n21 ), .ZN(\Check1_CheckInst_0_n23 ) );
  XNOR2_X1 \Check1_CheckInst_0_U26  ( .A(Red_ShiftRowsOutput[0]), .B(
        Red_SignaltoCheck[96]), .ZN(\Check1_CheckInst_0_n21 ) );
  XNOR2_X1 \Check1_CheckInst_0_U25  ( .A(Red_ShiftRowsOutput[3]), .B(
        Red_SignaltoCheck[99]), .ZN(\Check1_CheckInst_0_n22 ) );
  NAND2_X1 \Check1_CheckInst_0_U24  ( .A1(\Check1_CheckInst_0_n20 ), .A2(
        \Check1_CheckInst_0_n19 ), .ZN(\Check1_CheckInst_0_n24 ) );
  XNOR2_X1 \Check1_CheckInst_0_U23  ( .A(Red_Feedback[42]), .B(
        Red_SignaltoCheck[90]), .ZN(\Check1_CheckInst_0_n19 ) );
  XNOR2_X1 \Check1_CheckInst_0_U22  ( .A(Red_ShiftRowsOutput[6]), .B(
        Red_SignaltoCheck[102]), .ZN(\Check1_CheckInst_0_n20 ) );
  NOR2_X1 \Check1_CheckInst_0_U21  ( .A1(\Check1_CheckInst_0_n18 ), .A2(
        \Check1_CheckInst_0_n17 ), .ZN(\Check1_CheckInst_0_n26 ) );
  XOR2_X1 \Check1_CheckInst_0_U20  ( .A(Red_Feedback[45]), .B(
        Red_SignaltoCheck[93]), .Z(\Check1_CheckInst_0_n17 ) );
  XOR2_X1 \Check1_CheckInst_0_U19  ( .A(Red_Feedback[39]), .B(
        Red_SignaltoCheck[87]), .Z(\Check1_CheckInst_0_n18 ) );
  NAND2_X1 \Check1_CheckInst_0_U18  ( .A1(\Check1_CheckInst_0_n16 ), .A2(
        \Check1_CheckInst_0_n15 ), .ZN(\Check1_CheckInst_0_n28 ) );
  XNOR2_X1 \Check1_CheckInst_0_U17  ( .A(Red_Feedback[30]), .B(
        Red_SignaltoCheck[78]), .ZN(\Check1_CheckInst_0_n15 ) );
  XNOR2_X1 \Check1_CheckInst_0_U16  ( .A(Red_Feedback[33]), .B(
        Red_SignaltoCheck[81]), .ZN(\Check1_CheckInst_0_n16 ) );
  NAND2_X1 \Check1_CheckInst_0_U15  ( .A1(\Check1_CheckInst_0_n14 ), .A2(
        \Check1_CheckInst_0_n13 ), .ZN(\Check1_CheckInst_0_n94 ) );
  NOR2_X1 \Check1_CheckInst_0_U14  ( .A1(\Check1_CheckInst_0_n12 ), .A2(
        \Check1_CheckInst_0_n11 ), .ZN(\Check1_CheckInst_0_n13 ) );
  NAND2_X1 \Check1_CheckInst_0_U13  ( .A1(\Check1_CheckInst_0_n10 ), .A2(
        \Check1_CheckInst_0_n9 ), .ZN(\Check1_CheckInst_0_n11 ) );
  NOR2_X1 \Check1_CheckInst_0_U12  ( .A1(\Check1_CheckInst_0_n8 ), .A2(
        \Check1_CheckInst_0_n7 ), .ZN(\Check1_CheckInst_0_n9 ) );
  XOR2_X1 \Check1_CheckInst_0_U11  ( .A(Red_Feedback[24]), .B(
        Red_SignaltoCheck[72]), .Z(\Check1_CheckInst_0_n7 ) );
  XOR2_X1 \Check1_CheckInst_0_U10  ( .A(Red_Feedback[36]), .B(
        Red_SignaltoCheck[84]), .Z(\Check1_CheckInst_0_n8 ) );
  NOR2_X1 \Check1_CheckInst_0_U9  ( .A1(\Check1_CheckInst_0_n6 ), .A2(
        \Check1_CheckInst_0_n5 ), .ZN(\Check1_CheckInst_0_n10 ) );
  XOR2_X1 \Check1_CheckInst_0_U8  ( .A(Red_Feedback[27]), .B(
        Red_SignaltoCheck[75]), .Z(\Check1_CheckInst_0_n5 ) );
  XOR2_X1 \Check1_CheckInst_0_U7  ( .A(Red_Feedback[21]), .B(
        Red_SignaltoCheck[69]), .Z(\Check1_CheckInst_0_n6 ) );
  NAND2_X1 \Check1_CheckInst_0_U6  ( .A1(\Check1_CheckInst_0_n4 ), .A2(
        \Check1_CheckInst_0_n3 ), .ZN(\Check1_CheckInst_0_n12 ) );
  XNOR2_X1 \Check1_CheckInst_0_U5  ( .A(Red_ShiftRowsOutput[36]), .B(
        Red_SignaltoCheck[132]), .ZN(\Check1_CheckInst_0_n3 ) );
  XNOR2_X1 \Check1_CheckInst_0_U4  ( .A(Red_ShiftRowsOutput[39]), .B(
        Red_SignaltoCheck[135]), .ZN(\Check1_CheckInst_0_n4 ) );
  NOR2_X1 \Check1_CheckInst_0_U3  ( .A1(\Check1_CheckInst_0_n2 ), .A2(
        \Check1_CheckInst_0_n1 ), .ZN(\Check1_CheckInst_0_n14 ) );
  XOR2_X1 \Check1_CheckInst_0_U2  ( .A(Red_ShiftRowsOutput[30]), .B(
        Red_SignaltoCheck[126]), .Z(\Check1_CheckInst_0_n1 ) );
  XOR2_X1 \Check1_CheckInst_0_U1  ( .A(Red_ShiftRowsOutput[42]), .B(
        Red_SignaltoCheck[138]), .Z(\Check1_CheckInst_0_n2 ) );
  NOR2_X1 \Check1_CheckInst_1_U95  ( .A1(\Check1_CheckInst_1_n96 ), .A2(
        \Check1_CheckInst_1_n95 ), .ZN(Error[1]) );
  NAND2_X1 \Check1_CheckInst_1_U94  ( .A1(\Check1_CheckInst_1_n94 ), .A2(
        \Check1_CheckInst_1_n93 ), .ZN(\Check1_CheckInst_1_n95 ) );
  NOR2_X1 \Check1_CheckInst_1_U93  ( .A1(\Check1_CheckInst_1_n92 ), .A2(
        \Check1_CheckInst_1_n91 ), .ZN(\Check1_CheckInst_1_n93 ) );
  NAND2_X1 \Check1_CheckInst_1_U92  ( .A1(\Check1_CheckInst_1_n90 ), .A2(
        \Check1_CheckInst_1_n89 ), .ZN(\Check1_CheckInst_1_n91 ) );
  NOR2_X1 \Check1_CheckInst_1_U91  ( .A1(\Check1_CheckInst_1_n88 ), .A2(
        \Check1_CheckInst_1_n87 ), .ZN(\Check1_CheckInst_1_n89 ) );
  NAND2_X1 \Check1_CheckInst_1_U90  ( .A1(\Check1_CheckInst_1_n86 ), .A2(
        \Check1_CheckInst_1_n85 ), .ZN(\Check1_CheckInst_1_n87 ) );
  NOR2_X1 \Check1_CheckInst_1_U89  ( .A1(\Check1_CheckInst_1_n84 ), .A2(
        \Check1_CheckInst_1_n83 ), .ZN(\Check1_CheckInst_1_n85 ) );
  NAND2_X1 \Check1_CheckInst_1_U88  ( .A1(\Check1_CheckInst_1_n82 ), .A2(
        \Check1_CheckInst_1_n81 ), .ZN(\Check1_CheckInst_1_n83 ) );
  XNOR2_X1 \Check1_CheckInst_1_U87  ( .A(Red_ShiftRowsOutput[19]), .B(
        Red_SignaltoCheck[115]), .ZN(\Check1_CheckInst_1_n81 ) );
  XNOR2_X1 \Check1_CheckInst_1_U86  ( .A(Red_ShiftRowsOutput[22]), .B(
        Red_SignaltoCheck[118]), .ZN(\Check1_CheckInst_1_n82 ) );
  NAND2_X1 \Check1_CheckInst_1_U85  ( .A1(\Check1_CheckInst_1_n80 ), .A2(
        \Check1_CheckInst_1_n79 ), .ZN(\Check1_CheckInst_1_n84 ) );
  XNOR2_X1 \Check1_CheckInst_1_U84  ( .A(Red_ShiftRowsOutput[34]), .B(
        Red_SignaltoCheck[130]), .ZN(\Check1_CheckInst_1_n79 ) );
  XNOR2_X1 \Check1_CheckInst_1_U83  ( .A(Red_ShiftRowsOutput[28]), .B(
        Red_SignaltoCheck[124]), .ZN(\Check1_CheckInst_1_n80 ) );
  NOR2_X1 \Check1_CheckInst_1_U82  ( .A1(\Check1_CheckInst_1_n78 ), .A2(
        \Check1_CheckInst_1_n77 ), .ZN(\Check1_CheckInst_1_n86 ) );
  NAND2_X1 \Check1_CheckInst_1_U81  ( .A1(\Check1_CheckInst_1_n76 ), .A2(
        \Check1_CheckInst_1_n75 ), .ZN(\Check1_CheckInst_1_n77 ) );
  XNOR2_X1 \Check1_CheckInst_1_U80  ( .A(Red_ShiftRowsOutput[16]), .B(
        Red_SignaltoCheck[112]), .ZN(\Check1_CheckInst_1_n75 ) );
  XNOR2_X1 \Check1_CheckInst_1_U79  ( .A(Red_ShiftRowsOutput[10]), .B(
        Red_SignaltoCheck[106]), .ZN(\Check1_CheckInst_1_n76 ) );
  NAND2_X1 \Check1_CheckInst_1_U78  ( .A1(\Check1_CheckInst_1_n74 ), .A2(
        \Check1_CheckInst_1_n73 ), .ZN(\Check1_CheckInst_1_n78 ) );
  XNOR2_X1 \Check1_CheckInst_1_U77  ( .A(Red_ShiftRowsOutput[13]), .B(
        Red_SignaltoCheck[109]), .ZN(\Check1_CheckInst_1_n73 ) );
  XNOR2_X1 \Check1_CheckInst_1_U76  ( .A(Red_ShiftRowsOutput[25]), .B(
        Red_SignaltoCheck[121]), .ZN(\Check1_CheckInst_1_n74 ) );
  NAND2_X1 \Check1_CheckInst_1_U75  ( .A1(\Check1_CheckInst_1_n72 ), .A2(
        \Check1_CheckInst_1_n71 ), .ZN(\Check1_CheckInst_1_n88 ) );
  NOR2_X1 \Check1_CheckInst_1_U74  ( .A1(\Check1_CheckInst_1_n70 ), .A2(
        \Check1_CheckInst_1_n69 ), .ZN(\Check1_CheckInst_1_n71 ) );
  XOR2_X1 \Check1_CheckInst_1_U73  ( .A(Red_AddConstOutput[7]), .B(
        Red_SignaltoCheck[19]), .Z(\Check1_CheckInst_1_n69 ) );
  XOR2_X1 \Check1_CheckInst_1_U72  ( .A(Red_AddConstOutput[13]), .B(
        Red_SignaltoCheck[31]), .Z(\Check1_CheckInst_1_n70 ) );
  NOR2_X1 \Check1_CheckInst_1_U71  ( .A1(\Check1_CheckInst_1_n68 ), .A2(
        \Check1_CheckInst_1_n67 ), .ZN(\Check1_CheckInst_1_n72 ) );
  XOR2_X1 \Check1_CheckInst_1_U70  ( .A(Red_StateRegOutput[25]), .B(
        Red_SignaltoCheck[25]), .Z(\Check1_CheckInst_1_n67 ) );
  XOR2_X1 \Check1_CheckInst_1_U69  ( .A(Red_StateRegOutput[28]), .B(
        Red_SignaltoCheck[28]), .Z(\Check1_CheckInst_1_n68 ) );
  NOR2_X1 \Check1_CheckInst_1_U68  ( .A1(\Check1_CheckInst_1_n66 ), .A2(
        \Check1_CheckInst_1_n65 ), .ZN(\Check1_CheckInst_1_n90 ) );
  NAND2_X1 \Check1_CheckInst_1_U67  ( .A1(\Check1_CheckInst_1_n64 ), .A2(
        \Check1_CheckInst_1_n63 ), .ZN(\Check1_CheckInst_1_n65 ) );
  XNOR2_X1 \Check1_CheckInst_1_U66  ( .A(Red_AddConstOutput[1]), .B(
        Red_SignaltoCheck[7]), .ZN(\Check1_CheckInst_1_n63 ) );
  XNOR2_X1 \Check1_CheckInst_1_U65  ( .A(Red_AddConstOutput[4]), .B(
        Red_SignaltoCheck[10]), .ZN(\Check1_CheckInst_1_n64 ) );
  NAND2_X1 \Check1_CheckInst_1_U64  ( .A1(\Check1_CheckInst_1_n62 ), .A2(
        \Check1_CheckInst_1_n61 ), .ZN(\Check1_CheckInst_1_n66 ) );
  XNOR2_X1 \Check1_CheckInst_1_U63  ( .A(Red_AddConstOutput[10]), .B(
        Red_SignaltoCheck[22]), .ZN(\Check1_CheckInst_1_n61 ) );
  XNOR2_X1 \Check1_CheckInst_1_U62  ( .A(Red_StateRegOutput[16]), .B(
        Red_SignaltoCheck[16]), .ZN(\Check1_CheckInst_1_n62 ) );
  NAND2_X1 \Check1_CheckInst_1_U61  ( .A1(\Check1_CheckInst_1_n60 ), .A2(
        \Check1_CheckInst_1_n59 ), .ZN(\Check1_CheckInst_1_n92 ) );
  NOR2_X1 \Check1_CheckInst_1_U60  ( .A1(\Check1_CheckInst_1_n58 ), .A2(
        \Check1_CheckInst_1_n57 ), .ZN(\Check1_CheckInst_1_n59 ) );
  NAND2_X1 \Check1_CheckInst_1_U59  ( .A1(\Check1_CheckInst_1_n56 ), .A2(
        \Check1_CheckInst_1_n55 ), .ZN(\Check1_CheckInst_1_n57 ) );
  NOR2_X1 \Check1_CheckInst_1_U58  ( .A1(\Check1_CheckInst_1_n54 ), .A2(
        \Check1_CheckInst_1_n53 ), .ZN(\Check1_CheckInst_1_n55 ) );
  NAND2_X1 \Check1_CheckInst_1_U57  ( .A1(\Check1_CheckInst_1_n52 ), .A2(
        \Check1_CheckInst_1_n51 ), .ZN(\Check1_CheckInst_1_n53 ) );
  XNOR2_X1 \Check1_CheckInst_1_U56  ( .A(Red_ShiftRowsOutput[46]), .B(
        Red_SignaltoCheck[142]), .ZN(\Check1_CheckInst_1_n51 ) );
  XNOR2_X1 \Check1_CheckInst_1_U55  ( .A(Red_SignaltoCheck[4]), .B(
        Red_StateRegOutput[4]), .ZN(\Check1_CheckInst_1_n52 ) );
  NAND2_X1 \Check1_CheckInst_1_U54  ( .A1(\Check1_CheckInst_1_n50 ), .A2(
        \Check1_CheckInst_1_n49 ), .ZN(\Check1_CheckInst_1_n54 ) );
  XNOR2_X1 \Check1_CheckInst_1_U53  ( .A(Red_StateRegOutput[1]), .B(
        Red_SignaltoCheck[1]), .ZN(\Check1_CheckInst_1_n49 ) );
  XNOR2_X1 \Check1_CheckInst_1_U52  ( .A(Red_StateRegOutput[13]), .B(
        Red_SignaltoCheck[13]), .ZN(\Check1_CheckInst_1_n50 ) );
  NOR2_X1 \Check1_CheckInst_1_U51  ( .A1(\Check1_CheckInst_1_n48 ), .A2(
        \Check1_CheckInst_1_n47 ), .ZN(\Check1_CheckInst_1_n56 ) );
  NAND2_X1 \Check1_CheckInst_1_U50  ( .A1(\Check1_CheckInst_1_n46 ), .A2(
        \Check1_CheckInst_1_n45 ), .ZN(\Check1_CheckInst_1_n47 ) );
  XNOR2_X1 \Check1_CheckInst_1_U49  ( .A(Red_Feedback[7]), .B(
        Red_SignaltoCheck[55]), .ZN(\Check1_CheckInst_1_n45 ) );
  XNOR2_X1 \Check1_CheckInst_1_U48  ( .A(Red_Feedback[19]), .B(
        Red_SignaltoCheck[67]), .ZN(\Check1_CheckInst_1_n46 ) );
  NAND2_X1 \Check1_CheckInst_1_U47  ( .A1(\Check1_CheckInst_1_n44 ), .A2(
        \Check1_CheckInst_1_n43 ), .ZN(\Check1_CheckInst_1_n48 ) );
  XNOR2_X1 \Check1_CheckInst_1_U46  ( .A(Red_Feedback[13]), .B(
        Red_SignaltoCheck[61]), .ZN(\Check1_CheckInst_1_n43 ) );
  XNOR2_X1 \Check1_CheckInst_1_U45  ( .A(Red_Feedback[16]), .B(
        Red_SignaltoCheck[64]), .ZN(\Check1_CheckInst_1_n44 ) );
  NAND2_X1 \Check1_CheckInst_1_U44  ( .A1(\Check1_CheckInst_1_n42 ), .A2(
        \Check1_CheckInst_1_n41 ), .ZN(\Check1_CheckInst_1_n58 ) );
  NOR2_X1 \Check1_CheckInst_1_U43  ( .A1(\Check1_CheckInst_1_n40 ), .A2(
        \Check1_CheckInst_1_n39 ), .ZN(\Check1_CheckInst_1_n41 ) );
  XOR2_X1 \Check1_CheckInst_1_U42  ( .A(Red_AddConstOutput[19]), .B(
        Red_SignaltoCheck[43]), .Z(\Check1_CheckInst_1_n39 ) );
  XOR2_X1 \Check1_CheckInst_1_U41  ( .A(Red_AddConstOutput[22]), .B(
        Red_SignaltoCheck[46]), .Z(\Check1_CheckInst_1_n40 ) );
  NOR2_X1 \Check1_CheckInst_1_U40  ( .A1(\Check1_CheckInst_1_n38 ), .A2(
        \Check1_CheckInst_1_n37 ), .ZN(\Check1_CheckInst_1_n42 ) );
  XOR2_X1 \Check1_CheckInst_1_U39  ( .A(Red_Feedback[10]), .B(
        Red_SignaltoCheck[58]), .Z(\Check1_CheckInst_1_n37 ) );
  XOR2_X1 \Check1_CheckInst_1_U38  ( .A(Red_Feedback[4]), .B(
        Red_SignaltoCheck[52]), .Z(\Check1_CheckInst_1_n38 ) );
  NOR2_X1 \Check1_CheckInst_1_U37  ( .A1(\Check1_CheckInst_1_n36 ), .A2(
        \Check1_CheckInst_1_n35 ), .ZN(\Check1_CheckInst_1_n60 ) );
  NAND2_X1 \Check1_CheckInst_1_U36  ( .A1(\Check1_CheckInst_1_n34 ), .A2(
        \Check1_CheckInst_1_n33 ), .ZN(\Check1_CheckInst_1_n35 ) );
  XNOR2_X1 \Check1_CheckInst_1_U35  ( .A(Red_StateRegOutput[40]), .B(
        Red_SignaltoCheck[40]), .ZN(\Check1_CheckInst_1_n33 ) );
  XNOR2_X1 \Check1_CheckInst_1_U34  ( .A(Red_AddConstOutput[16]), .B(
        Red_SignaltoCheck[34]), .ZN(\Check1_CheckInst_1_n34 ) );
  NAND2_X1 \Check1_CheckInst_1_U33  ( .A1(\Check1_CheckInst_1_n32 ), .A2(
        \Check1_CheckInst_1_n31 ), .ZN(\Check1_CheckInst_1_n36 ) );
  XNOR2_X1 \Check1_CheckInst_1_U32  ( .A(Red_StateRegOutput[37]), .B(
        Red_SignaltoCheck[37]), .ZN(\Check1_CheckInst_1_n31 ) );
  XNOR2_X1 \Check1_CheckInst_1_U31  ( .A(Red_Feedback[1]), .B(
        Red_SignaltoCheck[49]), .ZN(\Check1_CheckInst_1_n32 ) );
  NOR2_X1 \Check1_CheckInst_1_U30  ( .A1(\Check1_CheckInst_1_n30 ), .A2(
        \Check1_CheckInst_1_n29 ), .ZN(\Check1_CheckInst_1_n94 ) );
  NAND2_X1 \Check1_CheckInst_1_U29  ( .A1(\Check1_CheckInst_1_n28 ), .A2(
        \Check1_CheckInst_1_n27 ), .ZN(\Check1_CheckInst_1_n29 ) );
  NOR2_X1 \Check1_CheckInst_1_U28  ( .A1(\Check1_CheckInst_1_n26 ), .A2(
        \Check1_CheckInst_1_n25 ), .ZN(\Check1_CheckInst_1_n27 ) );
  NAND2_X1 \Check1_CheckInst_1_U27  ( .A1(\Check1_CheckInst_1_n24 ), .A2(
        \Check1_CheckInst_1_n23 ), .ZN(\Check1_CheckInst_1_n25 ) );
  XNOR2_X1 \Check1_CheckInst_1_U26  ( .A(Red_ShiftRowsOutput[1]), .B(
        Red_SignaltoCheck[97]), .ZN(\Check1_CheckInst_1_n23 ) );
  XNOR2_X1 \Check1_CheckInst_1_U25  ( .A(Red_ShiftRowsOutput[4]), .B(
        Red_SignaltoCheck[100]), .ZN(\Check1_CheckInst_1_n24 ) );
  NAND2_X1 \Check1_CheckInst_1_U24  ( .A1(\Check1_CheckInst_1_n22 ), .A2(
        \Check1_CheckInst_1_n21 ), .ZN(\Check1_CheckInst_1_n26 ) );
  XNOR2_X1 \Check1_CheckInst_1_U23  ( .A(Red_Feedback[43]), .B(
        Red_SignaltoCheck[91]), .ZN(\Check1_CheckInst_1_n21 ) );
  XNOR2_X1 \Check1_CheckInst_1_U22  ( .A(Red_ShiftRowsOutput[7]), .B(
        Red_SignaltoCheck[103]), .ZN(\Check1_CheckInst_1_n22 ) );
  NOR2_X1 \Check1_CheckInst_1_U21  ( .A1(\Check1_CheckInst_1_n20 ), .A2(
        \Check1_CheckInst_1_n19 ), .ZN(\Check1_CheckInst_1_n28 ) );
  XOR2_X1 \Check1_CheckInst_1_U20  ( .A(Red_Feedback[46]), .B(
        Red_SignaltoCheck[94]), .Z(\Check1_CheckInst_1_n19 ) );
  XOR2_X1 \Check1_CheckInst_1_U19  ( .A(Red_Feedback[40]), .B(
        Red_SignaltoCheck[88]), .Z(\Check1_CheckInst_1_n20 ) );
  NAND2_X1 \Check1_CheckInst_1_U18  ( .A1(\Check1_CheckInst_1_n18 ), .A2(
        \Check1_CheckInst_1_n17 ), .ZN(\Check1_CheckInst_1_n30 ) );
  XNOR2_X1 \Check1_CheckInst_1_U17  ( .A(Red_Feedback[31]), .B(
        Red_SignaltoCheck[79]), .ZN(\Check1_CheckInst_1_n17 ) );
  XNOR2_X1 \Check1_CheckInst_1_U16  ( .A(Red_Feedback[34]), .B(
        Red_SignaltoCheck[82]), .ZN(\Check1_CheckInst_1_n18 ) );
  NAND2_X1 \Check1_CheckInst_1_U15  ( .A1(\Check1_CheckInst_1_n16 ), .A2(
        \Check1_CheckInst_1_n15 ), .ZN(\Check1_CheckInst_1_n96 ) );
  NOR2_X1 \Check1_CheckInst_1_U14  ( .A1(\Check1_CheckInst_1_n14 ), .A2(
        \Check1_CheckInst_1_n13 ), .ZN(\Check1_CheckInst_1_n15 ) );
  NAND2_X1 \Check1_CheckInst_1_U13  ( .A1(\Check1_CheckInst_1_n12 ), .A2(
        \Check1_CheckInst_1_n11 ), .ZN(\Check1_CheckInst_1_n13 ) );
  NOR2_X1 \Check1_CheckInst_1_U12  ( .A1(\Check1_CheckInst_1_n10 ), .A2(
        \Check1_CheckInst_1_n9 ), .ZN(\Check1_CheckInst_1_n11 ) );
  XOR2_X1 \Check1_CheckInst_1_U11  ( .A(Red_Feedback[25]), .B(
        Red_SignaltoCheck[73]), .Z(\Check1_CheckInst_1_n9 ) );
  XOR2_X1 \Check1_CheckInst_1_U10  ( .A(Red_Feedback[37]), .B(
        Red_SignaltoCheck[85]), .Z(\Check1_CheckInst_1_n10 ) );
  NOR2_X1 \Check1_CheckInst_1_U9  ( .A1(\Check1_CheckInst_1_n8 ), .A2(
        \Check1_CheckInst_1_n7 ), .ZN(\Check1_CheckInst_1_n12 ) );
  XOR2_X1 \Check1_CheckInst_1_U8  ( .A(Red_Feedback[28]), .B(
        Red_SignaltoCheck[76]), .Z(\Check1_CheckInst_1_n7 ) );
  XOR2_X1 \Check1_CheckInst_1_U7  ( .A(Red_Feedback[22]), .B(
        Red_SignaltoCheck[70]), .Z(\Check1_CheckInst_1_n8 ) );
  NAND2_X1 \Check1_CheckInst_1_U6  ( .A1(\Check1_CheckInst_1_n6 ), .A2(
        \Check1_CheckInst_1_n5 ), .ZN(\Check1_CheckInst_1_n14 ) );
  XNOR2_X1 \Check1_CheckInst_1_U5  ( .A(Red_ShiftRowsOutput[37]), .B(
        Red_SignaltoCheck[133]), .ZN(\Check1_CheckInst_1_n5 ) );
  XNOR2_X1 \Check1_CheckInst_1_U4  ( .A(Red_ShiftRowsOutput[40]), .B(
        Red_SignaltoCheck[136]), .ZN(\Check1_CheckInst_1_n6 ) );
  NOR2_X1 \Check1_CheckInst_1_U3  ( .A1(\Check1_CheckInst_1_n4 ), .A2(
        \Check1_CheckInst_1_n3 ), .ZN(\Check1_CheckInst_1_n16 ) );
  XOR2_X1 \Check1_CheckInst_1_U2  ( .A(Red_ShiftRowsOutput[31]), .B(
        Red_SignaltoCheck[127]), .Z(\Check1_CheckInst_1_n3 ) );
  XOR2_X1 \Check1_CheckInst_1_U1  ( .A(Red_ShiftRowsOutput[43]), .B(
        Red_SignaltoCheck[139]), .Z(\Check1_CheckInst_1_n4 ) );
  NOR2_X1 \Check1_CheckInst_2_U95  ( .A1(\Check1_CheckInst_2_n96 ), .A2(
        \Check1_CheckInst_2_n95 ), .ZN(Error[2]) );
  NAND2_X1 \Check1_CheckInst_2_U94  ( .A1(\Check1_CheckInst_2_n94 ), .A2(
        \Check1_CheckInst_2_n93 ), .ZN(\Check1_CheckInst_2_n95 ) );
  NOR2_X1 \Check1_CheckInst_2_U93  ( .A1(\Check1_CheckInst_2_n92 ), .A2(
        \Check1_CheckInst_2_n91 ), .ZN(\Check1_CheckInst_2_n93 ) );
  NAND2_X1 \Check1_CheckInst_2_U92  ( .A1(\Check1_CheckInst_2_n90 ), .A2(
        \Check1_CheckInst_2_n89 ), .ZN(\Check1_CheckInst_2_n91 ) );
  NOR2_X1 \Check1_CheckInst_2_U91  ( .A1(\Check1_CheckInst_2_n88 ), .A2(
        \Check1_CheckInst_2_n87 ), .ZN(\Check1_CheckInst_2_n89 ) );
  NAND2_X1 \Check1_CheckInst_2_U90  ( .A1(\Check1_CheckInst_2_n86 ), .A2(
        \Check1_CheckInst_2_n85 ), .ZN(\Check1_CheckInst_2_n87 ) );
  NOR2_X1 \Check1_CheckInst_2_U89  ( .A1(\Check1_CheckInst_2_n84 ), .A2(
        \Check1_CheckInst_2_n83 ), .ZN(\Check1_CheckInst_2_n85 ) );
  NAND2_X1 \Check1_CheckInst_2_U88  ( .A1(\Check1_CheckInst_2_n82 ), .A2(
        \Check1_CheckInst_2_n81 ), .ZN(\Check1_CheckInst_2_n83 ) );
  XNOR2_X1 \Check1_CheckInst_2_U87  ( .A(Red_ShiftRowsOutput[20]), .B(
        Red_SignaltoCheck[116]), .ZN(\Check1_CheckInst_2_n81 ) );
  XNOR2_X1 \Check1_CheckInst_2_U86  ( .A(Red_ShiftRowsOutput[23]), .B(
        Red_SignaltoCheck[119]), .ZN(\Check1_CheckInst_2_n82 ) );
  NAND2_X1 \Check1_CheckInst_2_U85  ( .A1(\Check1_CheckInst_2_n80 ), .A2(
        \Check1_CheckInst_2_n79 ), .ZN(\Check1_CheckInst_2_n84 ) );
  XNOR2_X1 \Check1_CheckInst_2_U84  ( .A(Red_ShiftRowsOutput[35]), .B(
        Red_SignaltoCheck[131]), .ZN(\Check1_CheckInst_2_n79 ) );
  XNOR2_X1 \Check1_CheckInst_2_U83  ( .A(Red_ShiftRowsOutput[29]), .B(
        Red_SignaltoCheck[125]), .ZN(\Check1_CheckInst_2_n80 ) );
  NOR2_X1 \Check1_CheckInst_2_U82  ( .A1(\Check1_CheckInst_2_n78 ), .A2(
        \Check1_CheckInst_2_n77 ), .ZN(\Check1_CheckInst_2_n86 ) );
  NAND2_X1 \Check1_CheckInst_2_U81  ( .A1(\Check1_CheckInst_2_n76 ), .A2(
        \Check1_CheckInst_2_n75 ), .ZN(\Check1_CheckInst_2_n77 ) );
  XNOR2_X1 \Check1_CheckInst_2_U80  ( .A(Red_ShiftRowsOutput[17]), .B(
        Red_SignaltoCheck[113]), .ZN(\Check1_CheckInst_2_n75 ) );
  XNOR2_X1 \Check1_CheckInst_2_U79  ( .A(Red_ShiftRowsOutput[11]), .B(
        Red_SignaltoCheck[107]), .ZN(\Check1_CheckInst_2_n76 ) );
  NAND2_X1 \Check1_CheckInst_2_U78  ( .A1(\Check1_CheckInst_2_n74 ), .A2(
        \Check1_CheckInst_2_n73 ), .ZN(\Check1_CheckInst_2_n78 ) );
  XNOR2_X1 \Check1_CheckInst_2_U77  ( .A(Red_ShiftRowsOutput[14]), .B(
        Red_SignaltoCheck[110]), .ZN(\Check1_CheckInst_2_n73 ) );
  XNOR2_X1 \Check1_CheckInst_2_U76  ( .A(Red_ShiftRowsOutput[26]), .B(
        Red_SignaltoCheck[122]), .ZN(\Check1_CheckInst_2_n74 ) );
  NAND2_X1 \Check1_CheckInst_2_U75  ( .A1(\Check1_CheckInst_2_n72 ), .A2(
        \Check1_CheckInst_2_n71 ), .ZN(\Check1_CheckInst_2_n88 ) );
  NOR2_X1 \Check1_CheckInst_2_U74  ( .A1(\Check1_CheckInst_2_n70 ), .A2(
        \Check1_CheckInst_2_n69 ), .ZN(\Check1_CheckInst_2_n71 ) );
  XOR2_X1 \Check1_CheckInst_2_U73  ( .A(Red_AddConstOutput[8]), .B(
        Red_SignaltoCheck[20]), .Z(\Check1_CheckInst_2_n69 ) );
  XOR2_X1 \Check1_CheckInst_2_U72  ( .A(Red_AddConstOutput[14]), .B(
        Red_SignaltoCheck[32]), .Z(\Check1_CheckInst_2_n70 ) );
  NOR2_X1 \Check1_CheckInst_2_U71  ( .A1(\Check1_CheckInst_2_n68 ), .A2(
        \Check1_CheckInst_2_n67 ), .ZN(\Check1_CheckInst_2_n72 ) );
  XOR2_X1 \Check1_CheckInst_2_U70  ( .A(Red_StateRegOutput[26]), .B(
        Red_SignaltoCheck[26]), .Z(\Check1_CheckInst_2_n67 ) );
  XOR2_X1 \Check1_CheckInst_2_U69  ( .A(Red_StateRegOutput[29]), .B(
        Red_SignaltoCheck[29]), .Z(\Check1_CheckInst_2_n68 ) );
  NOR2_X1 \Check1_CheckInst_2_U68  ( .A1(\Check1_CheckInst_2_n66 ), .A2(
        \Check1_CheckInst_2_n65 ), .ZN(\Check1_CheckInst_2_n90 ) );
  NAND2_X1 \Check1_CheckInst_2_U67  ( .A1(\Check1_CheckInst_2_n64 ), .A2(
        \Check1_CheckInst_2_n63 ), .ZN(\Check1_CheckInst_2_n65 ) );
  XNOR2_X1 \Check1_CheckInst_2_U66  ( .A(Red_AddConstOutput[2]), .B(
        Red_SignaltoCheck[8]), .ZN(\Check1_CheckInst_2_n63 ) );
  XNOR2_X1 \Check1_CheckInst_2_U65  ( .A(Red_AddConstOutput[5]), .B(
        Red_SignaltoCheck[11]), .ZN(\Check1_CheckInst_2_n64 ) );
  NAND2_X1 \Check1_CheckInst_2_U64  ( .A1(\Check1_CheckInst_2_n62 ), .A2(
        \Check1_CheckInst_2_n61 ), .ZN(\Check1_CheckInst_2_n66 ) );
  XNOR2_X1 \Check1_CheckInst_2_U63  ( .A(Red_AddConstOutput[11]), .B(
        Red_SignaltoCheck[23]), .ZN(\Check1_CheckInst_2_n61 ) );
  XNOR2_X1 \Check1_CheckInst_2_U62  ( .A(Red_StateRegOutput[17]), .B(
        Red_SignaltoCheck[17]), .ZN(\Check1_CheckInst_2_n62 ) );
  NAND2_X1 \Check1_CheckInst_2_U61  ( .A1(\Check1_CheckInst_2_n60 ), .A2(
        \Check1_CheckInst_2_n59 ), .ZN(\Check1_CheckInst_2_n92 ) );
  NOR2_X1 \Check1_CheckInst_2_U60  ( .A1(\Check1_CheckInst_2_n58 ), .A2(
        \Check1_CheckInst_2_n57 ), .ZN(\Check1_CheckInst_2_n59 ) );
  NAND2_X1 \Check1_CheckInst_2_U59  ( .A1(\Check1_CheckInst_2_n56 ), .A2(
        \Check1_CheckInst_2_n55 ), .ZN(\Check1_CheckInst_2_n57 ) );
  NOR2_X1 \Check1_CheckInst_2_U58  ( .A1(\Check1_CheckInst_2_n54 ), .A2(
        \Check1_CheckInst_2_n53 ), .ZN(\Check1_CheckInst_2_n55 ) );
  NAND2_X1 \Check1_CheckInst_2_U57  ( .A1(\Check1_CheckInst_2_n52 ), .A2(
        \Check1_CheckInst_2_n51 ), .ZN(\Check1_CheckInst_2_n53 ) );
  XNOR2_X1 \Check1_CheckInst_2_U56  ( .A(Red_ShiftRowsOutput[47]), .B(
        Red_SignaltoCheck[143]), .ZN(\Check1_CheckInst_2_n51 ) );
  XNOR2_X1 \Check1_CheckInst_2_U55  ( .A(Red_SignaltoCheck[5]), .B(
        Red_StateRegOutput[5]), .ZN(\Check1_CheckInst_2_n52 ) );
  NAND2_X1 \Check1_CheckInst_2_U54  ( .A1(\Check1_CheckInst_2_n50 ), .A2(
        \Check1_CheckInst_2_n49 ), .ZN(\Check1_CheckInst_2_n54 ) );
  XNOR2_X1 \Check1_CheckInst_2_U53  ( .A(Red_StateRegOutput[2]), .B(
        Red_SignaltoCheck[2]), .ZN(\Check1_CheckInst_2_n49 ) );
  XNOR2_X1 \Check1_CheckInst_2_U52  ( .A(Red_StateRegOutput[14]), .B(
        Red_SignaltoCheck[14]), .ZN(\Check1_CheckInst_2_n50 ) );
  NOR2_X1 \Check1_CheckInst_2_U51  ( .A1(\Check1_CheckInst_2_n48 ), .A2(
        \Check1_CheckInst_2_n47 ), .ZN(\Check1_CheckInst_2_n56 ) );
  NAND2_X1 \Check1_CheckInst_2_U50  ( .A1(\Check1_CheckInst_2_n46 ), .A2(
        \Check1_CheckInst_2_n45 ), .ZN(\Check1_CheckInst_2_n47 ) );
  XNOR2_X1 \Check1_CheckInst_2_U49  ( .A(Red_Feedback[8]), .B(
        Red_SignaltoCheck[56]), .ZN(\Check1_CheckInst_2_n45 ) );
  XNOR2_X1 \Check1_CheckInst_2_U48  ( .A(Red_Feedback[20]), .B(
        Red_SignaltoCheck[68]), .ZN(\Check1_CheckInst_2_n46 ) );
  NAND2_X1 \Check1_CheckInst_2_U47  ( .A1(\Check1_CheckInst_2_n44 ), .A2(
        \Check1_CheckInst_2_n43 ), .ZN(\Check1_CheckInst_2_n48 ) );
  XNOR2_X1 \Check1_CheckInst_2_U46  ( .A(Red_Feedback[14]), .B(
        Red_SignaltoCheck[62]), .ZN(\Check1_CheckInst_2_n43 ) );
  XNOR2_X1 \Check1_CheckInst_2_U45  ( .A(Red_Feedback[17]), .B(
        Red_SignaltoCheck[65]), .ZN(\Check1_CheckInst_2_n44 ) );
  NAND2_X1 \Check1_CheckInst_2_U44  ( .A1(\Check1_CheckInst_2_n42 ), .A2(
        \Check1_CheckInst_2_n41 ), .ZN(\Check1_CheckInst_2_n58 ) );
  NOR2_X1 \Check1_CheckInst_2_U43  ( .A1(\Check1_CheckInst_2_n40 ), .A2(
        \Check1_CheckInst_2_n39 ), .ZN(\Check1_CheckInst_2_n41 ) );
  XOR2_X1 \Check1_CheckInst_2_U42  ( .A(Red_AddConstOutput[20]), .B(
        Red_SignaltoCheck[44]), .Z(\Check1_CheckInst_2_n39 ) );
  XOR2_X1 \Check1_CheckInst_2_U41  ( .A(Red_AddConstOutput[23]), .B(
        Red_SignaltoCheck[47]), .Z(\Check1_CheckInst_2_n40 ) );
  NOR2_X1 \Check1_CheckInst_2_U40  ( .A1(\Check1_CheckInst_2_n38 ), .A2(
        \Check1_CheckInst_2_n37 ), .ZN(\Check1_CheckInst_2_n42 ) );
  XOR2_X1 \Check1_CheckInst_2_U39  ( .A(Red_Feedback[11]), .B(
        Red_SignaltoCheck[59]), .Z(\Check1_CheckInst_2_n37 ) );
  XOR2_X1 \Check1_CheckInst_2_U38  ( .A(Red_Feedback[5]), .B(
        Red_SignaltoCheck[53]), .Z(\Check1_CheckInst_2_n38 ) );
  NOR2_X1 \Check1_CheckInst_2_U37  ( .A1(\Check1_CheckInst_2_n36 ), .A2(
        \Check1_CheckInst_2_n35 ), .ZN(\Check1_CheckInst_2_n60 ) );
  NAND2_X1 \Check1_CheckInst_2_U36  ( .A1(\Check1_CheckInst_2_n34 ), .A2(
        \Check1_CheckInst_2_n33 ), .ZN(\Check1_CheckInst_2_n35 ) );
  XNOR2_X1 \Check1_CheckInst_2_U35  ( .A(Red_StateRegOutput[41]), .B(
        Red_SignaltoCheck[41]), .ZN(\Check1_CheckInst_2_n33 ) );
  XNOR2_X1 \Check1_CheckInst_2_U34  ( .A(Red_AddConstOutput[17]), .B(
        Red_SignaltoCheck[35]), .ZN(\Check1_CheckInst_2_n34 ) );
  NAND2_X1 \Check1_CheckInst_2_U33  ( .A1(\Check1_CheckInst_2_n32 ), .A2(
        \Check1_CheckInst_2_n31 ), .ZN(\Check1_CheckInst_2_n36 ) );
  XNOR2_X1 \Check1_CheckInst_2_U32  ( .A(Red_StateRegOutput[38]), .B(
        Red_SignaltoCheck[38]), .ZN(\Check1_CheckInst_2_n31 ) );
  XNOR2_X1 \Check1_CheckInst_2_U31  ( .A(Red_Feedback[2]), .B(
        Red_SignaltoCheck[50]), .ZN(\Check1_CheckInst_2_n32 ) );
  NOR2_X1 \Check1_CheckInst_2_U30  ( .A1(\Check1_CheckInst_2_n30 ), .A2(
        \Check1_CheckInst_2_n29 ), .ZN(\Check1_CheckInst_2_n94 ) );
  NAND2_X1 \Check1_CheckInst_2_U29  ( .A1(\Check1_CheckInst_2_n28 ), .A2(
        \Check1_CheckInst_2_n27 ), .ZN(\Check1_CheckInst_2_n29 ) );
  NOR2_X1 \Check1_CheckInst_2_U28  ( .A1(\Check1_CheckInst_2_n26 ), .A2(
        \Check1_CheckInst_2_n25 ), .ZN(\Check1_CheckInst_2_n27 ) );
  NAND2_X1 \Check1_CheckInst_2_U27  ( .A1(\Check1_CheckInst_2_n24 ), .A2(
        \Check1_CheckInst_2_n23 ), .ZN(\Check1_CheckInst_2_n25 ) );
  XNOR2_X1 \Check1_CheckInst_2_U26  ( .A(Red_ShiftRowsOutput[2]), .B(
        Red_SignaltoCheck[98]), .ZN(\Check1_CheckInst_2_n23 ) );
  XNOR2_X1 \Check1_CheckInst_2_U25  ( .A(Red_ShiftRowsOutput[5]), .B(
        Red_SignaltoCheck[101]), .ZN(\Check1_CheckInst_2_n24 ) );
  NAND2_X1 \Check1_CheckInst_2_U24  ( .A1(\Check1_CheckInst_2_n22 ), .A2(
        \Check1_CheckInst_2_n21 ), .ZN(\Check1_CheckInst_2_n26 ) );
  XNOR2_X1 \Check1_CheckInst_2_U23  ( .A(Red_Feedback[44]), .B(
        Red_SignaltoCheck[92]), .ZN(\Check1_CheckInst_2_n21 ) );
  XNOR2_X1 \Check1_CheckInst_2_U22  ( .A(Red_ShiftRowsOutput[8]), .B(
        Red_SignaltoCheck[104]), .ZN(\Check1_CheckInst_2_n22 ) );
  NOR2_X1 \Check1_CheckInst_2_U21  ( .A1(\Check1_CheckInst_2_n20 ), .A2(
        \Check1_CheckInst_2_n19 ), .ZN(\Check1_CheckInst_2_n28 ) );
  XOR2_X1 \Check1_CheckInst_2_U20  ( .A(Red_Feedback[47]), .B(
        Red_SignaltoCheck[95]), .Z(\Check1_CheckInst_2_n19 ) );
  XOR2_X1 \Check1_CheckInst_2_U19  ( .A(Red_Feedback[41]), .B(
        Red_SignaltoCheck[89]), .Z(\Check1_CheckInst_2_n20 ) );
  NAND2_X1 \Check1_CheckInst_2_U18  ( .A1(\Check1_CheckInst_2_n18 ), .A2(
        \Check1_CheckInst_2_n17 ), .ZN(\Check1_CheckInst_2_n30 ) );
  XNOR2_X1 \Check1_CheckInst_2_U17  ( .A(Red_Feedback[32]), .B(
        Red_SignaltoCheck[80]), .ZN(\Check1_CheckInst_2_n17 ) );
  XNOR2_X1 \Check1_CheckInst_2_U16  ( .A(Red_Feedback[35]), .B(
        Red_SignaltoCheck[83]), .ZN(\Check1_CheckInst_2_n18 ) );
  NAND2_X1 \Check1_CheckInst_2_U15  ( .A1(\Check1_CheckInst_2_n16 ), .A2(
        \Check1_CheckInst_2_n15 ), .ZN(\Check1_CheckInst_2_n96 ) );
  NOR2_X1 \Check1_CheckInst_2_U14  ( .A1(\Check1_CheckInst_2_n14 ), .A2(
        \Check1_CheckInst_2_n13 ), .ZN(\Check1_CheckInst_2_n15 ) );
  NAND2_X1 \Check1_CheckInst_2_U13  ( .A1(\Check1_CheckInst_2_n12 ), .A2(
        \Check1_CheckInst_2_n11 ), .ZN(\Check1_CheckInst_2_n13 ) );
  NOR2_X1 \Check1_CheckInst_2_U12  ( .A1(\Check1_CheckInst_2_n10 ), .A2(
        \Check1_CheckInst_2_n9 ), .ZN(\Check1_CheckInst_2_n11 ) );
  XOR2_X1 \Check1_CheckInst_2_U11  ( .A(Red_Feedback[26]), .B(
        Red_SignaltoCheck[74]), .Z(\Check1_CheckInst_2_n9 ) );
  XOR2_X1 \Check1_CheckInst_2_U10  ( .A(Red_Feedback[38]), .B(
        Red_SignaltoCheck[86]), .Z(\Check1_CheckInst_2_n10 ) );
  NOR2_X1 \Check1_CheckInst_2_U9  ( .A1(\Check1_CheckInst_2_n8 ), .A2(
        \Check1_CheckInst_2_n7 ), .ZN(\Check1_CheckInst_2_n12 ) );
  XOR2_X1 \Check1_CheckInst_2_U8  ( .A(Red_Feedback[29]), .B(
        Red_SignaltoCheck[77]), .Z(\Check1_CheckInst_2_n7 ) );
  XOR2_X1 \Check1_CheckInst_2_U7  ( .A(Red_Feedback[23]), .B(
        Red_SignaltoCheck[71]), .Z(\Check1_CheckInst_2_n8 ) );
  NAND2_X1 \Check1_CheckInst_2_U6  ( .A1(\Check1_CheckInst_2_n6 ), .A2(
        \Check1_CheckInst_2_n5 ), .ZN(\Check1_CheckInst_2_n14 ) );
  XNOR2_X1 \Check1_CheckInst_2_U5  ( .A(Red_ShiftRowsOutput[38]), .B(
        Red_SignaltoCheck[134]), .ZN(\Check1_CheckInst_2_n5 ) );
  XNOR2_X1 \Check1_CheckInst_2_U4  ( .A(Red_ShiftRowsOutput[41]), .B(
        Red_SignaltoCheck[137]), .ZN(\Check1_CheckInst_2_n6 ) );
  NOR2_X1 \Check1_CheckInst_2_U3  ( .A1(\Check1_CheckInst_2_n4 ), .A2(
        \Check1_CheckInst_2_n3 ), .ZN(\Check1_CheckInst_2_n16 ) );
  XOR2_X1 \Check1_CheckInst_2_U2  ( .A(Red_ShiftRowsOutput[32]), .B(
        Red_SignaltoCheck[128]), .Z(\Check1_CheckInst_2_n3 ) );
  XOR2_X1 \Check1_CheckInst_2_U1  ( .A(Red_ShiftRowsOutput[44]), .B(
        Red_SignaltoCheck[140]), .Z(\Check1_CheckInst_2_n4 ) );
endmodule

