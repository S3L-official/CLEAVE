module Cipher ( clk, rst, EncDec, Input, Key, Output, ErrorFlag );
  input [63:0] Input;
  input [63:0] Key;
  output [63:0] Output;
  (* FIRMER="clock" *)input clk, rst, EncDec;
  output ErrorFlag;
  wire   n8, n9, \MCInst_XOR_r0_Inst_0_n3 , \MCInst_XOR_r0_Inst_1_n3 ,
         \MCInst_XOR_r0_Inst_2_n3 , \MCInst_XOR_r0_Inst_3_n3 ,
         \MCInst_XOR_r0_Inst_4_n3 , \MCInst_XOR_r0_Inst_5_n3 ,
         \MCInst_XOR_r0_Inst_6_n3 , \MCInst_XOR_r0_Inst_7_n3 ,
         \MCInst_XOR_r0_Inst_8_n3 , \MCInst_XOR_r0_Inst_9_n3 ,
         \MCInst_XOR_r0_Inst_10_n3 , \MCInst_XOR_r0_Inst_11_n3 ,
         \MCInst_XOR_r0_Inst_12_n3 , \MCInst_XOR_r0_Inst_13_n3 ,
         \MCInst_XOR_r0_Inst_14_n3 , \MCInst_XOR_r0_Inst_15_n3 ,
         \SubCellInst_LFInst_0_LFInst_0_n11 ,
         \SubCellInst_LFInst_0_LFInst_0_n10 ,
         \SubCellInst_LFInst_0_LFInst_0_n9 ,
         \SubCellInst_LFInst_0_LFInst_0_n8 ,
         \SubCellInst_LFInst_0_LFInst_0_n7 ,
         \SubCellInst_LFInst_0_LFInst_1_n6 ,
         \SubCellInst_LFInst_0_LFInst_1_n5 ,
         \SubCellInst_LFInst_0_LFInst_1_n4 ,
         \SubCellInst_LFInst_0_LFInst_2_n11 ,
         \SubCellInst_LFInst_0_LFInst_2_n10 ,
         \SubCellInst_LFInst_0_LFInst_2_n9 ,
         \SubCellInst_LFInst_0_LFInst_2_n8 ,
         \SubCellInst_LFInst_0_LFInst_2_n7 ,
         \SubCellInst_LFInst_0_LFInst_3_n6 ,
         \SubCellInst_LFInst_0_LFInst_3_n5 ,
         \SubCellInst_LFInst_0_LFInst_3_n4 ,
         \SubCellInst_LFInst_1_LFInst_0_n11 ,
         \SubCellInst_LFInst_1_LFInst_0_n10 ,
         \SubCellInst_LFInst_1_LFInst_0_n9 ,
         \SubCellInst_LFInst_1_LFInst_0_n8 ,
         \SubCellInst_LFInst_1_LFInst_0_n7 ,
         \SubCellInst_LFInst_1_LFInst_1_n6 ,
         \SubCellInst_LFInst_1_LFInst_1_n5 ,
         \SubCellInst_LFInst_1_LFInst_1_n4 ,
         \SubCellInst_LFInst_1_LFInst_2_n11 ,
         \SubCellInst_LFInst_1_LFInst_2_n10 ,
         \SubCellInst_LFInst_1_LFInst_2_n9 ,
         \SubCellInst_LFInst_1_LFInst_2_n8 ,
         \SubCellInst_LFInst_1_LFInst_2_n7 ,
         \SubCellInst_LFInst_1_LFInst_3_n6 ,
         \SubCellInst_LFInst_1_LFInst_3_n5 ,
         \SubCellInst_LFInst_1_LFInst_3_n4 ,
         \SubCellInst_LFInst_2_LFInst_0_n11 ,
         \SubCellInst_LFInst_2_LFInst_0_n10 ,
         \SubCellInst_LFInst_2_LFInst_0_n9 ,
         \SubCellInst_LFInst_2_LFInst_0_n8 ,
         \SubCellInst_LFInst_2_LFInst_0_n7 ,
         \SubCellInst_LFInst_2_LFInst_1_n6 ,
         \SubCellInst_LFInst_2_LFInst_1_n5 ,
         \SubCellInst_LFInst_2_LFInst_1_n4 ,
         \SubCellInst_LFInst_2_LFInst_2_n11 ,
         \SubCellInst_LFInst_2_LFInst_2_n10 ,
         \SubCellInst_LFInst_2_LFInst_2_n9 ,
         \SubCellInst_LFInst_2_LFInst_2_n8 ,
         \SubCellInst_LFInst_2_LFInst_2_n7 ,
         \SubCellInst_LFInst_2_LFInst_3_n6 ,
         \SubCellInst_LFInst_2_LFInst_3_n5 ,
         \SubCellInst_LFInst_2_LFInst_3_n4 ,
         \SubCellInst_LFInst_3_LFInst_0_n11 ,
         \SubCellInst_LFInst_3_LFInst_0_n10 ,
         \SubCellInst_LFInst_3_LFInst_0_n9 ,
         \SubCellInst_LFInst_3_LFInst_0_n8 ,
         \SubCellInst_LFInst_3_LFInst_0_n7 ,
         \SubCellInst_LFInst_3_LFInst_1_n6 ,
         \SubCellInst_LFInst_3_LFInst_1_n5 ,
         \SubCellInst_LFInst_3_LFInst_1_n4 ,
         \SubCellInst_LFInst_3_LFInst_2_n11 ,
         \SubCellInst_LFInst_3_LFInst_2_n10 ,
         \SubCellInst_LFInst_3_LFInst_2_n9 ,
         \SubCellInst_LFInst_3_LFInst_2_n8 ,
         \SubCellInst_LFInst_3_LFInst_2_n7 ,
         \SubCellInst_LFInst_3_LFInst_3_n6 ,
         \SubCellInst_LFInst_3_LFInst_3_n5 ,
         \SubCellInst_LFInst_3_LFInst_3_n4 ,
         \SubCellInst_LFInst_4_LFInst_0_n11 ,
         \SubCellInst_LFInst_4_LFInst_0_n10 ,
         \SubCellInst_LFInst_4_LFInst_0_n9 ,
         \SubCellInst_LFInst_4_LFInst_0_n8 ,
         \SubCellInst_LFInst_4_LFInst_0_n7 ,
         \SubCellInst_LFInst_4_LFInst_1_n6 ,
         \SubCellInst_LFInst_4_LFInst_1_n5 ,
         \SubCellInst_LFInst_4_LFInst_1_n4 ,
         \SubCellInst_LFInst_4_LFInst_2_n11 ,
         \SubCellInst_LFInst_4_LFInst_2_n10 ,
         \SubCellInst_LFInst_4_LFInst_2_n9 ,
         \SubCellInst_LFInst_4_LFInst_2_n8 ,
         \SubCellInst_LFInst_4_LFInst_2_n7 ,
         \SubCellInst_LFInst_4_LFInst_3_n6 ,
         \SubCellInst_LFInst_4_LFInst_3_n5 ,
         \SubCellInst_LFInst_4_LFInst_3_n4 ,
         \SubCellInst_LFInst_5_LFInst_0_n11 ,
         \SubCellInst_LFInst_5_LFInst_0_n10 ,
         \SubCellInst_LFInst_5_LFInst_0_n9 ,
         \SubCellInst_LFInst_5_LFInst_0_n8 ,
         \SubCellInst_LFInst_5_LFInst_0_n7 ,
         \SubCellInst_LFInst_5_LFInst_1_n6 ,
         \SubCellInst_LFInst_5_LFInst_1_n5 ,
         \SubCellInst_LFInst_5_LFInst_1_n4 ,
         \SubCellInst_LFInst_5_LFInst_2_n11 ,
         \SubCellInst_LFInst_5_LFInst_2_n10 ,
         \SubCellInst_LFInst_5_LFInst_2_n9 ,
         \SubCellInst_LFInst_5_LFInst_2_n8 ,
         \SubCellInst_LFInst_5_LFInst_2_n7 ,
         \SubCellInst_LFInst_5_LFInst_3_n6 ,
         \SubCellInst_LFInst_5_LFInst_3_n5 ,
         \SubCellInst_LFInst_5_LFInst_3_n4 ,
         \SubCellInst_LFInst_6_LFInst_0_n11 ,
         \SubCellInst_LFInst_6_LFInst_0_n10 ,
         \SubCellInst_LFInst_6_LFInst_0_n9 ,
         \SubCellInst_LFInst_6_LFInst_0_n8 ,
         \SubCellInst_LFInst_6_LFInst_0_n7 ,
         \SubCellInst_LFInst_6_LFInst_1_n6 ,
         \SubCellInst_LFInst_6_LFInst_1_n5 ,
         \SubCellInst_LFInst_6_LFInst_1_n4 ,
         \SubCellInst_LFInst_6_LFInst_2_n11 ,
         \SubCellInst_LFInst_6_LFInst_2_n10 ,
         \SubCellInst_LFInst_6_LFInst_2_n9 ,
         \SubCellInst_LFInst_6_LFInst_2_n8 ,
         \SubCellInst_LFInst_6_LFInst_2_n7 ,
         \SubCellInst_LFInst_6_LFInst_3_n6 ,
         \SubCellInst_LFInst_6_LFInst_3_n5 ,
         \SubCellInst_LFInst_6_LFInst_3_n4 ,
         \SubCellInst_LFInst_7_LFInst_0_n11 ,
         \SubCellInst_LFInst_7_LFInst_0_n10 ,
         \SubCellInst_LFInst_7_LFInst_0_n9 ,
         \SubCellInst_LFInst_7_LFInst_0_n8 ,
         \SubCellInst_LFInst_7_LFInst_0_n7 ,
         \SubCellInst_LFInst_7_LFInst_1_n6 ,
         \SubCellInst_LFInst_7_LFInst_1_n5 ,
         \SubCellInst_LFInst_7_LFInst_1_n4 ,
         \SubCellInst_LFInst_7_LFInst_2_n11 ,
         \SubCellInst_LFInst_7_LFInst_2_n10 ,
         \SubCellInst_LFInst_7_LFInst_2_n9 ,
         \SubCellInst_LFInst_7_LFInst_2_n8 ,
         \SubCellInst_LFInst_7_LFInst_2_n7 ,
         \SubCellInst_LFInst_7_LFInst_3_n6 ,
         \SubCellInst_LFInst_7_LFInst_3_n5 ,
         \SubCellInst_LFInst_7_LFInst_3_n4 ,
         \SubCellInst_LFInst_8_LFInst_0_n11 ,
         \SubCellInst_LFInst_8_LFInst_0_n10 ,
         \SubCellInst_LFInst_8_LFInst_0_n9 ,
         \SubCellInst_LFInst_8_LFInst_0_n8 ,
         \SubCellInst_LFInst_8_LFInst_0_n7 ,
         \SubCellInst_LFInst_8_LFInst_1_n6 ,
         \SubCellInst_LFInst_8_LFInst_1_n5 ,
         \SubCellInst_LFInst_8_LFInst_1_n4 ,
         \SubCellInst_LFInst_8_LFInst_2_n11 ,
         \SubCellInst_LFInst_8_LFInst_2_n10 ,
         \SubCellInst_LFInst_8_LFInst_2_n9 ,
         \SubCellInst_LFInst_8_LFInst_2_n8 ,
         \SubCellInst_LFInst_8_LFInst_2_n7 ,
         \SubCellInst_LFInst_8_LFInst_3_n6 ,
         \SubCellInst_LFInst_8_LFInst_3_n5 ,
         \SubCellInst_LFInst_8_LFInst_3_n4 ,
         \SubCellInst_LFInst_9_LFInst_0_n11 ,
         \SubCellInst_LFInst_9_LFInst_0_n10 ,
         \SubCellInst_LFInst_9_LFInst_0_n9 ,
         \SubCellInst_LFInst_9_LFInst_0_n8 ,
         \SubCellInst_LFInst_9_LFInst_0_n7 ,
         \SubCellInst_LFInst_9_LFInst_1_n6 ,
         \SubCellInst_LFInst_9_LFInst_1_n5 ,
         \SubCellInst_LFInst_9_LFInst_1_n4 ,
         \SubCellInst_LFInst_9_LFInst_2_n11 ,
         \SubCellInst_LFInst_9_LFInst_2_n10 ,
         \SubCellInst_LFInst_9_LFInst_2_n9 ,
         \SubCellInst_LFInst_9_LFInst_2_n8 ,
         \SubCellInst_LFInst_9_LFInst_2_n7 ,
         \SubCellInst_LFInst_9_LFInst_3_n6 ,
         \SubCellInst_LFInst_9_LFInst_3_n5 ,
         \SubCellInst_LFInst_9_LFInst_3_n4 ,
         \SubCellInst_LFInst_10_LFInst_0_n11 ,
         \SubCellInst_LFInst_10_LFInst_0_n10 ,
         \SubCellInst_LFInst_10_LFInst_0_n9 ,
         \SubCellInst_LFInst_10_LFInst_0_n8 ,
         \SubCellInst_LFInst_10_LFInst_0_n7 ,
         \SubCellInst_LFInst_10_LFInst_1_n6 ,
         \SubCellInst_LFInst_10_LFInst_1_n5 ,
         \SubCellInst_LFInst_10_LFInst_1_n4 ,
         \SubCellInst_LFInst_10_LFInst_2_n11 ,
         \SubCellInst_LFInst_10_LFInst_2_n10 ,
         \SubCellInst_LFInst_10_LFInst_2_n9 ,
         \SubCellInst_LFInst_10_LFInst_2_n8 ,
         \SubCellInst_LFInst_10_LFInst_2_n7 ,
         \SubCellInst_LFInst_10_LFInst_3_n6 ,
         \SubCellInst_LFInst_10_LFInst_3_n5 ,
         \SubCellInst_LFInst_10_LFInst_3_n4 ,
         \SubCellInst_LFInst_11_LFInst_0_n11 ,
         \SubCellInst_LFInst_11_LFInst_0_n10 ,
         \SubCellInst_LFInst_11_LFInst_0_n9 ,
         \SubCellInst_LFInst_11_LFInst_0_n8 ,
         \SubCellInst_LFInst_11_LFInst_0_n7 ,
         \SubCellInst_LFInst_11_LFInst_1_n6 ,
         \SubCellInst_LFInst_11_LFInst_1_n5 ,
         \SubCellInst_LFInst_11_LFInst_1_n4 ,
         \SubCellInst_LFInst_11_LFInst_2_n11 ,
         \SubCellInst_LFInst_11_LFInst_2_n10 ,
         \SubCellInst_LFInst_11_LFInst_2_n9 ,
         \SubCellInst_LFInst_11_LFInst_2_n8 ,
         \SubCellInst_LFInst_11_LFInst_2_n7 ,
         \SubCellInst_LFInst_11_LFInst_3_n6 ,
         \SubCellInst_LFInst_11_LFInst_3_n5 ,
         \SubCellInst_LFInst_11_LFInst_3_n4 ,
         \SubCellInst_LFInst_12_LFInst_0_n11 ,
         \SubCellInst_LFInst_12_LFInst_0_n10 ,
         \SubCellInst_LFInst_12_LFInst_0_n9 ,
         \SubCellInst_LFInst_12_LFInst_0_n8 ,
         \SubCellInst_LFInst_12_LFInst_0_n7 ,
         \SubCellInst_LFInst_12_LFInst_1_n6 ,
         \SubCellInst_LFInst_12_LFInst_1_n5 ,
         \SubCellInst_LFInst_12_LFInst_1_n4 ,
         \SubCellInst_LFInst_12_LFInst_2_n11 ,
         \SubCellInst_LFInst_12_LFInst_2_n10 ,
         \SubCellInst_LFInst_12_LFInst_2_n9 ,
         \SubCellInst_LFInst_12_LFInst_2_n8 ,
         \SubCellInst_LFInst_12_LFInst_2_n7 ,
         \SubCellInst_LFInst_12_LFInst_3_n6 ,
         \SubCellInst_LFInst_12_LFInst_3_n5 ,
         \SubCellInst_LFInst_12_LFInst_3_n4 ,
         \SubCellInst_LFInst_13_LFInst_0_n11 ,
         \SubCellInst_LFInst_13_LFInst_0_n10 ,
         \SubCellInst_LFInst_13_LFInst_0_n9 ,
         \SubCellInst_LFInst_13_LFInst_0_n8 ,
         \SubCellInst_LFInst_13_LFInst_0_n7 ,
         \SubCellInst_LFInst_13_LFInst_1_n6 ,
         \SubCellInst_LFInst_13_LFInst_1_n5 ,
         \SubCellInst_LFInst_13_LFInst_1_n4 ,
         \SubCellInst_LFInst_13_LFInst_2_n11 ,
         \SubCellInst_LFInst_13_LFInst_2_n10 ,
         \SubCellInst_LFInst_13_LFInst_2_n9 ,
         \SubCellInst_LFInst_13_LFInst_2_n8 ,
         \SubCellInst_LFInst_13_LFInst_2_n7 ,
         \SubCellInst_LFInst_13_LFInst_3_n6 ,
         \SubCellInst_LFInst_13_LFInst_3_n5 ,
         \SubCellInst_LFInst_13_LFInst_3_n4 ,
         \SubCellInst_LFInst_14_LFInst_0_n11 ,
         \SubCellInst_LFInst_14_LFInst_0_n10 ,
         \SubCellInst_LFInst_14_LFInst_0_n9 ,
         \SubCellInst_LFInst_14_LFInst_0_n8 ,
         \SubCellInst_LFInst_14_LFInst_0_n7 ,
         \SubCellInst_LFInst_14_LFInst_1_n6 ,
         \SubCellInst_LFInst_14_LFInst_1_n5 ,
         \SubCellInst_LFInst_14_LFInst_1_n4 ,
         \SubCellInst_LFInst_14_LFInst_2_n11 ,
         \SubCellInst_LFInst_14_LFInst_2_n10 ,
         \SubCellInst_LFInst_14_LFInst_2_n9 ,
         \SubCellInst_LFInst_14_LFInst_2_n8 ,
         \SubCellInst_LFInst_14_LFInst_2_n7 ,
         \SubCellInst_LFInst_14_LFInst_3_n6 ,
         \SubCellInst_LFInst_14_LFInst_3_n5 ,
         \SubCellInst_LFInst_14_LFInst_3_n4 ,
         \SubCellInst_LFInst_15_LFInst_0_n11 ,
         \SubCellInst_LFInst_15_LFInst_0_n10 ,
         \SubCellInst_LFInst_15_LFInst_0_n9 ,
         \SubCellInst_LFInst_15_LFInst_0_n8 ,
         \SubCellInst_LFInst_15_LFInst_0_n7 ,
         \SubCellInst_LFInst_15_LFInst_1_n6 ,
         \SubCellInst_LFInst_15_LFInst_1_n5 ,
         \SubCellInst_LFInst_15_LFInst_1_n4 ,
         \SubCellInst_LFInst_15_LFInst_2_n11 ,
         \SubCellInst_LFInst_15_LFInst_2_n10 ,
         \SubCellInst_LFInst_15_LFInst_2_n9 ,
         \SubCellInst_LFInst_15_LFInst_2_n8 ,
         \SubCellInst_LFInst_15_LFInst_2_n7 ,
         \SubCellInst_LFInst_15_LFInst_3_n6 ,
         \SubCellInst_LFInst_15_LFInst_3_n5 ,
         \SubCellInst_LFInst_15_LFInst_3_n4 ,
         \Red_PlaintextInst_LFInst_0_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_0_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_0_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_0_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_1_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_1_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_1_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_1_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_2_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_2_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_2_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_2_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_3_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_3_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_3_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_3_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_4_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_4_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_4_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_4_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_5_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_5_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_5_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_5_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_6_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_6_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_6_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_6_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_7_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_7_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_7_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_7_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_8_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_8_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_8_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_8_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_9_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_9_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_9_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_9_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_10_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_10_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_10_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_10_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_11_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_11_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_11_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_11_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_12_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_12_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_12_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_12_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_13_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_13_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_13_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_13_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_14_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_14_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_14_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_14_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_15_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_15_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_15_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_15_LFInst_3_n2 ,
         \Red_MCInst_XOR_r0_Inst_0_n3 , \Red_MCInst_XOR_r0_Inst_1_n3 ,
         \Red_MCInst_XOR_r0_Inst_2_n3 , \Red_MCInst_XOR_r0_Inst_3_n3 ,
         \Red_MCInst_XOR_r0_Inst_4_n3 , \Red_MCInst_XOR_r0_Inst_5_n3 ,
         \Red_MCInst_XOR_r0_Inst_6_n3 , \Red_MCInst_XOR_r0_Inst_7_n3 ,
         \Red_MCInst_XOR_r0_Inst_8_n3 , \Red_MCInst_XOR_r0_Inst_9_n3 ,
         \Red_MCInst_XOR_r0_Inst_10_n3 , \Red_MCInst_XOR_r0_Inst_11_n3 ,
         \Red_MCInst_XOR_r0_Inst_12_n3 , \Red_MCInst_XOR_r0_Inst_13_n3 ,
         \Red_MCInst_XOR_r0_Inst_14_n3 , \Red_MCInst_XOR_r0_Inst_15_n3 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_0_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_0_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_0_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_0_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_0_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_0_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_0_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_0_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_1_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_1_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_1_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_1_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_1_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_1_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_1_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_1_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_2_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_2_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_2_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_2_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_2_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_2_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_2_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_2_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_3_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_3_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_3_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_3_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_3_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_3_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_3_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_3_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_4_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_4_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_4_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_4_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_4_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_4_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_4_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_4_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_5_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_5_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_5_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_5_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_5_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_5_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_5_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_5_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_6_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_6_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_6_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_6_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_6_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_6_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_6_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_6_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_7_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_7_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_7_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_7_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_7_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_7_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_7_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_7_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_8_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_8_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_8_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_8_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_8_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_8_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_8_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_8_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_9_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_9_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_9_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_9_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_9_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_9_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_9_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_9_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_10_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_10_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_10_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_10_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_10_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_10_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_10_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_10_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_11_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_11_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_11_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_11_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_11_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_11_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_11_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_11_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_12_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_12_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_12_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_12_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_12_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_12_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_12_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_12_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_13_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_13_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_13_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_13_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_13_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_13_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_13_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_13_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_14_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_14_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_14_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_14_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_14_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_14_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_14_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_14_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_15_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_15_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_15_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_15_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_15_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_15_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_15_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_15_LFInst_3_n6 ,
         \Red_K0Inst_LFInst_0_LFInst_0_n2 , \Red_K0Inst_LFInst_0_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_0_LFInst_2_n2 , \Red_K0Inst_LFInst_0_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_1_LFInst_0_n2 , \Red_K0Inst_LFInst_1_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_1_LFInst_2_n2 , \Red_K0Inst_LFInst_1_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_2_LFInst_0_n2 , \Red_K0Inst_LFInst_2_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_2_LFInst_2_n2 , \Red_K0Inst_LFInst_2_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_3_LFInst_0_n2 , \Red_K0Inst_LFInst_3_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_3_LFInst_2_n2 , \Red_K0Inst_LFInst_3_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_4_LFInst_0_n2 , \Red_K0Inst_LFInst_4_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_4_LFInst_2_n2 , \Red_K0Inst_LFInst_4_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_5_LFInst_0_n2 , \Red_K0Inst_LFInst_5_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_5_LFInst_2_n2 , \Red_K0Inst_LFInst_5_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_6_LFInst_0_n2 , \Red_K0Inst_LFInst_6_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_6_LFInst_2_n2 , \Red_K0Inst_LFInst_6_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_7_LFInst_0_n2 , \Red_K0Inst_LFInst_7_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_7_LFInst_2_n2 , \Red_K0Inst_LFInst_7_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_8_LFInst_0_n2 , \Red_K0Inst_LFInst_8_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_8_LFInst_2_n2 , \Red_K0Inst_LFInst_8_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_9_LFInst_0_n2 , \Red_K0Inst_LFInst_9_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_9_LFInst_2_n2 , \Red_K0Inst_LFInst_9_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_10_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_10_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_10_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_10_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_11_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_11_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_11_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_11_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_12_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_12_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_12_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_12_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_13_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_13_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_13_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_13_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_14_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_14_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_14_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_14_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_15_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_15_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_15_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_15_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_0_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_0_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_0_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_0_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_1_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_1_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_1_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_1_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_2_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_2_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_2_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_2_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_3_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_3_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_3_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_3_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_4_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_4_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_4_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_4_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_5_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_5_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_5_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_5_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_6_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_6_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_6_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_6_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_7_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_7_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_7_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_7_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_8_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_8_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_8_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_8_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_9_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_9_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_9_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_9_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_10_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_10_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_10_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_10_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_11_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_11_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_11_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_11_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_12_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_12_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_12_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_12_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_13_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_13_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_13_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_13_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_14_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_14_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_14_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_14_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_15_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_15_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_15_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_15_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_16_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_16_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_16_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_16_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_17_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_17_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_17_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_17_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_18_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_18_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_18_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_18_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_19_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_19_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_19_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_19_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_20_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_20_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_20_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_20_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_21_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_21_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_21_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_21_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_22_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_22_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_22_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_22_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_23_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_23_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_23_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_23_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_24_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_24_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_24_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_24_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_25_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_25_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_25_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_25_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_26_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_26_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_26_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_26_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_27_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_27_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_27_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_27_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_28_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_28_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_28_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_28_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_29_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_29_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_29_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_29_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_30_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_30_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_30_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_30_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_31_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_31_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_31_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_31_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_32_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_32_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_32_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_32_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_33_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_33_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_33_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_33_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_34_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_34_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_34_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_34_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_35_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_35_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_35_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_35_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_36_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_36_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_36_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_36_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_37_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_37_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_37_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_37_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_38_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_38_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_38_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_38_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_39_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_39_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_39_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_39_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_40_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_40_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_40_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_40_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_41_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_41_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_41_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_41_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_42_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_42_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_42_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_42_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_43_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_43_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_43_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_43_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_44_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_44_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_44_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_44_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_45_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_45_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_45_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_45_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_46_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_46_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_46_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_46_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_47_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_47_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_47_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_47_LFInst_3_n2 , \Check1_CheckInst_0_n94 ,
         \Check1_CheckInst_0_n93 , \Check1_CheckInst_0_n92 ,
         \Check1_CheckInst_0_n91 , \Check1_CheckInst_0_n90 ,
         \Check1_CheckInst_0_n89 , \Check1_CheckInst_0_n88 ,
         \Check1_CheckInst_0_n87 , \Check1_CheckInst_0_n86 ,
         \Check1_CheckInst_0_n85 , \Check1_CheckInst_0_n84 ,
         \Check1_CheckInst_0_n83 , \Check1_CheckInst_0_n82 ,
         \Check1_CheckInst_0_n81 , \Check1_CheckInst_0_n80 ,
         \Check1_CheckInst_0_n79 , \Check1_CheckInst_0_n78 ,
         \Check1_CheckInst_0_n77 , \Check1_CheckInst_0_n76 ,
         \Check1_CheckInst_0_n75 , \Check1_CheckInst_0_n74 ,
         \Check1_CheckInst_0_n73 , \Check1_CheckInst_0_n72 ,
         \Check1_CheckInst_0_n71 , \Check1_CheckInst_0_n70 ,
         \Check1_CheckInst_0_n69 , \Check1_CheckInst_0_n68 ,
         \Check1_CheckInst_0_n67 , \Check1_CheckInst_0_n66 ,
         \Check1_CheckInst_0_n65 , \Check1_CheckInst_0_n64 ,
         \Check1_CheckInst_0_n63 , \Check1_CheckInst_0_n62 ,
         \Check1_CheckInst_0_n61 , \Check1_CheckInst_0_n60 ,
         \Check1_CheckInst_0_n59 , \Check1_CheckInst_0_n58 ,
         \Check1_CheckInst_0_n57 , \Check1_CheckInst_0_n56 ,
         \Check1_CheckInst_0_n55 , \Check1_CheckInst_0_n54 ,
         \Check1_CheckInst_0_n53 , \Check1_CheckInst_0_n52 ,
         \Check1_CheckInst_0_n51 , \Check1_CheckInst_0_n50 ,
         \Check1_CheckInst_0_n49 , \Check1_CheckInst_0_n48 ,
         \Check1_CheckInst_0_n47 , \Check1_CheckInst_0_n46 ,
         \Check1_CheckInst_0_n45 , \Check1_CheckInst_0_n44 ,
         \Check1_CheckInst_0_n43 , \Check1_CheckInst_0_n42 ,
         \Check1_CheckInst_0_n41 , \Check1_CheckInst_0_n40 ,
         \Check1_CheckInst_0_n39 , \Check1_CheckInst_0_n38 ,
         \Check1_CheckInst_0_n37 , \Check1_CheckInst_0_n36 ,
         \Check1_CheckInst_0_n35 , \Check1_CheckInst_0_n34 ,
         \Check1_CheckInst_0_n33 , \Check1_CheckInst_0_n32 ,
         \Check1_CheckInst_0_n31 , \Check1_CheckInst_0_n30 ,
         \Check1_CheckInst_0_n29 , \Check1_CheckInst_0_n28 ,
         \Check1_CheckInst_0_n27 , \Check1_CheckInst_0_n26 ,
         \Check1_CheckInst_0_n25 , \Check1_CheckInst_0_n24 ,
         \Check1_CheckInst_0_n23 , \Check1_CheckInst_0_n22 ,
         \Check1_CheckInst_0_n21 , \Check1_CheckInst_0_n20 ,
         \Check1_CheckInst_0_n19 , \Check1_CheckInst_0_n18 ,
         \Check1_CheckInst_0_n17 , \Check1_CheckInst_0_n16 ,
         \Check1_CheckInst_0_n15 , \Check1_CheckInst_0_n14 ,
         \Check1_CheckInst_0_n13 , \Check1_CheckInst_0_n12 ,
         \Check1_CheckInst_0_n11 , \Check1_CheckInst_0_n10 ,
         \Check1_CheckInst_0_n9 , \Check1_CheckInst_0_n8 ,
         \Check1_CheckInst_0_n7 , \Check1_CheckInst_0_n6 ,
         \Check1_CheckInst_0_n5 , \Check1_CheckInst_0_n4 ,
         \Check1_CheckInst_0_n3 , \Check1_CheckInst_0_n2 ,
         \Check1_CheckInst_0_n1 , \Check1_CheckInst_1_n96 ,
         \Check1_CheckInst_1_n95 , \Check1_CheckInst_1_n94 ,
         \Check1_CheckInst_1_n93 , \Check1_CheckInst_1_n92 ,
         \Check1_CheckInst_1_n91 , \Check1_CheckInst_1_n90 ,
         \Check1_CheckInst_1_n89 , \Check1_CheckInst_1_n88 ,
         \Check1_CheckInst_1_n87 , \Check1_CheckInst_1_n86 ,
         \Check1_CheckInst_1_n85 , \Check1_CheckInst_1_n84 ,
         \Check1_CheckInst_1_n83 , \Check1_CheckInst_1_n82 ,
         \Check1_CheckInst_1_n81 , \Check1_CheckInst_1_n80 ,
         \Check1_CheckInst_1_n79 , \Check1_CheckInst_1_n78 ,
         \Check1_CheckInst_1_n77 , \Check1_CheckInst_1_n76 ,
         \Check1_CheckInst_1_n75 , \Check1_CheckInst_1_n74 ,
         \Check1_CheckInst_1_n73 , \Check1_CheckInst_1_n72 ,
         \Check1_CheckInst_1_n71 , \Check1_CheckInst_1_n70 ,
         \Check1_CheckInst_1_n69 , \Check1_CheckInst_1_n68 ,
         \Check1_CheckInst_1_n67 , \Check1_CheckInst_1_n66 ,
         \Check1_CheckInst_1_n65 , \Check1_CheckInst_1_n64 ,
         \Check1_CheckInst_1_n63 , \Check1_CheckInst_1_n62 ,
         \Check1_CheckInst_1_n61 , \Check1_CheckInst_1_n60 ,
         \Check1_CheckInst_1_n59 , \Check1_CheckInst_1_n58 ,
         \Check1_CheckInst_1_n57 , \Check1_CheckInst_1_n56 ,
         \Check1_CheckInst_1_n55 , \Check1_CheckInst_1_n54 ,
         \Check1_CheckInst_1_n53 , \Check1_CheckInst_1_n52 ,
         \Check1_CheckInst_1_n51 , \Check1_CheckInst_1_n50 ,
         \Check1_CheckInst_1_n49 , \Check1_CheckInst_1_n48 ,
         \Check1_CheckInst_1_n47 , \Check1_CheckInst_1_n46 ,
         \Check1_CheckInst_1_n45 , \Check1_CheckInst_1_n44 ,
         \Check1_CheckInst_1_n43 , \Check1_CheckInst_1_n42 ,
         \Check1_CheckInst_1_n41 , \Check1_CheckInst_1_n40 ,
         \Check1_CheckInst_1_n39 , \Check1_CheckInst_1_n38 ,
         \Check1_CheckInst_1_n37 , \Check1_CheckInst_1_n36 ,
         \Check1_CheckInst_1_n35 , \Check1_CheckInst_1_n34 ,
         \Check1_CheckInst_1_n33 , \Check1_CheckInst_1_n32 ,
         \Check1_CheckInst_1_n31 , \Check1_CheckInst_1_n30 ,
         \Check1_CheckInst_1_n29 , \Check1_CheckInst_1_n28 ,
         \Check1_CheckInst_1_n27 , \Check1_CheckInst_1_n26 ,
         \Check1_CheckInst_1_n25 , \Check1_CheckInst_1_n24 ,
         \Check1_CheckInst_1_n23 , \Check1_CheckInst_1_n22 ,
         \Check1_CheckInst_1_n21 , \Check1_CheckInst_1_n20 ,
         \Check1_CheckInst_1_n19 , \Check1_CheckInst_1_n18 ,
         \Check1_CheckInst_1_n17 , \Check1_CheckInst_1_n16 ,
         \Check1_CheckInst_1_n15 , \Check1_CheckInst_1_n14 ,
         \Check1_CheckInst_1_n13 , \Check1_CheckInst_1_n12 ,
         \Check1_CheckInst_1_n11 , \Check1_CheckInst_1_n10 ,
         \Check1_CheckInst_1_n9 , \Check1_CheckInst_1_n8 ,
         \Check1_CheckInst_1_n7 , \Check1_CheckInst_1_n6 ,
         \Check1_CheckInst_1_n5 , \Check1_CheckInst_1_n4 ,
         \Check1_CheckInst_1_n3 , \Check1_CheckInst_2_n96 ,
         \Check1_CheckInst_2_n95 , \Check1_CheckInst_2_n94 ,
         \Check1_CheckInst_2_n93 , \Check1_CheckInst_2_n92 ,
         \Check1_CheckInst_2_n91 , \Check1_CheckInst_2_n90 ,
         \Check1_CheckInst_2_n89 , \Check1_CheckInst_2_n88 ,
         \Check1_CheckInst_2_n87 , \Check1_CheckInst_2_n86 ,
         \Check1_CheckInst_2_n85 , \Check1_CheckInst_2_n84 ,
         \Check1_CheckInst_2_n83 , \Check1_CheckInst_2_n82 ,
         \Check1_CheckInst_2_n81 , \Check1_CheckInst_2_n80 ,
         \Check1_CheckInst_2_n79 , \Check1_CheckInst_2_n78 ,
         \Check1_CheckInst_2_n77 , \Check1_CheckInst_2_n76 ,
         \Check1_CheckInst_2_n75 , \Check1_CheckInst_2_n74 ,
         \Check1_CheckInst_2_n73 , \Check1_CheckInst_2_n72 ,
         \Check1_CheckInst_2_n71 , \Check1_CheckInst_2_n70 ,
         \Check1_CheckInst_2_n69 , \Check1_CheckInst_2_n68 ,
         \Check1_CheckInst_2_n67 , \Check1_CheckInst_2_n66 ,
         \Check1_CheckInst_2_n65 , \Check1_CheckInst_2_n64 ,
         \Check1_CheckInst_2_n63 , \Check1_CheckInst_2_n62 ,
         \Check1_CheckInst_2_n61 , \Check1_CheckInst_2_n60 ,
         \Check1_CheckInst_2_n59 , \Check1_CheckInst_2_n58 ,
         \Check1_CheckInst_2_n57 , \Check1_CheckInst_2_n56 ,
         \Check1_CheckInst_2_n55 , \Check1_CheckInst_2_n54 ,
         \Check1_CheckInst_2_n53 , \Check1_CheckInst_2_n52 ,
         \Check1_CheckInst_2_n51 , \Check1_CheckInst_2_n50 ,
         \Check1_CheckInst_2_n49 , \Check1_CheckInst_2_n48 ,
         \Check1_CheckInst_2_n47 , \Check1_CheckInst_2_n46 ,
         \Check1_CheckInst_2_n45 , \Check1_CheckInst_2_n44 ,
         \Check1_CheckInst_2_n43 , \Check1_CheckInst_2_n42 ,
         \Check1_CheckInst_2_n41 , \Check1_CheckInst_2_n40 ,
         \Check1_CheckInst_2_n39 , \Check1_CheckInst_2_n38 ,
         \Check1_CheckInst_2_n37 , \Check1_CheckInst_2_n36 ,
         \Check1_CheckInst_2_n35 , \Check1_CheckInst_2_n34 ,
         \Check1_CheckInst_2_n33 , \Check1_CheckInst_2_n32 ,
         \Check1_CheckInst_2_n31 , \Check1_CheckInst_2_n30 ,
         \Check1_CheckInst_2_n29 , \Check1_CheckInst_2_n28 ,
         \Check1_CheckInst_2_n27 , \Check1_CheckInst_2_n26 ,
         \Check1_CheckInst_2_n25 , \Check1_CheckInst_2_n24 ,
         \Check1_CheckInst_2_n23 , \Check1_CheckInst_2_n22 ,
         \Check1_CheckInst_2_n21 , \Check1_CheckInst_2_n20 ,
         \Check1_CheckInst_2_n19 , \Check1_CheckInst_2_n18 ,
         \Check1_CheckInst_2_n17 , \Check1_CheckInst_2_n16 ,
         \Check1_CheckInst_2_n15 , \Check1_CheckInst_2_n14 ,
         \Check1_CheckInst_2_n13 , \Check1_CheckInst_2_n12 ,
         \Check1_CheckInst_2_n11 , \Check1_CheckInst_2_n10 ,
         \Check1_CheckInst_2_n9 , \Check1_CheckInst_2_n8 ,
         \Check1_CheckInst_2_n7 , \Check1_CheckInst_2_n6 ,
         \Check1_CheckInst_2_n5 , \Check1_CheckInst_2_n4 ,
         \Check1_CheckInst_2_n3 , \Check1_CheckInst_3_n96 ,
         \Check1_CheckInst_3_n95 , \Check1_CheckInst_3_n94 ,
         \Check1_CheckInst_3_n93 , \Check1_CheckInst_3_n92 ,
         \Check1_CheckInst_3_n91 , \Check1_CheckInst_3_n90 ,
         \Check1_CheckInst_3_n89 , \Check1_CheckInst_3_n88 ,
         \Check1_CheckInst_3_n87 , \Check1_CheckInst_3_n86 ,
         \Check1_CheckInst_3_n85 , \Check1_CheckInst_3_n84 ,
         \Check1_CheckInst_3_n83 , \Check1_CheckInst_3_n82 ,
         \Check1_CheckInst_3_n81 , \Check1_CheckInst_3_n80 ,
         \Check1_CheckInst_3_n79 , \Check1_CheckInst_3_n78 ,
         \Check1_CheckInst_3_n77 , \Check1_CheckInst_3_n76 ,
         \Check1_CheckInst_3_n75 , \Check1_CheckInst_3_n74 ,
         \Check1_CheckInst_3_n73 , \Check1_CheckInst_3_n72 ,
         \Check1_CheckInst_3_n71 , \Check1_CheckInst_3_n70 ,
         \Check1_CheckInst_3_n69 , \Check1_CheckInst_3_n68 ,
         \Check1_CheckInst_3_n67 , \Check1_CheckInst_3_n66 ,
         \Check1_CheckInst_3_n65 , \Check1_CheckInst_3_n64 ,
         \Check1_CheckInst_3_n63 , \Check1_CheckInst_3_n62 ,
         \Check1_CheckInst_3_n61 , \Check1_CheckInst_3_n60 ,
         \Check1_CheckInst_3_n59 , \Check1_CheckInst_3_n58 ,
         \Check1_CheckInst_3_n57 , \Check1_CheckInst_3_n56 ,
         \Check1_CheckInst_3_n55 , \Check1_CheckInst_3_n54 ,
         \Check1_CheckInst_3_n53 , \Check1_CheckInst_3_n52 ,
         \Check1_CheckInst_3_n51 , \Check1_CheckInst_3_n50 ,
         \Check1_CheckInst_3_n49 , \Check1_CheckInst_3_n48 ,
         \Check1_CheckInst_3_n47 , \Check1_CheckInst_3_n46 ,
         \Check1_CheckInst_3_n45 , \Check1_CheckInst_3_n44 ,
         \Check1_CheckInst_3_n43 , \Check1_CheckInst_3_n42 ,
         \Check1_CheckInst_3_n41 , \Check1_CheckInst_3_n40 ,
         \Check1_CheckInst_3_n39 , \Check1_CheckInst_3_n38 ,
         \Check1_CheckInst_3_n37 , \Check1_CheckInst_3_n36 ,
         \Check1_CheckInst_3_n35 , \Check1_CheckInst_3_n34 ,
         \Check1_CheckInst_3_n33 , \Check1_CheckInst_3_n32 ,
         \Check1_CheckInst_3_n31 , \Check1_CheckInst_3_n30 ,
         \Check1_CheckInst_3_n29 , \Check1_CheckInst_3_n28 ,
         \Check1_CheckInst_3_n27 , \Check1_CheckInst_3_n26 ,
         \Check1_CheckInst_3_n25 , \Check1_CheckInst_3_n24 ,
         \Check1_CheckInst_3_n23 , \Check1_CheckInst_3_n22 ,
         \Check1_CheckInst_3_n21 , \Check1_CheckInst_3_n20 ,
         \Check1_CheckInst_3_n19 , \Check1_CheckInst_3_n18 ,
         \Check1_CheckInst_3_n17 , \Check1_CheckInst_3_n16 ,
         \Check1_CheckInst_3_n15 , \Check1_CheckInst_3_n14 ,
         \Check1_CheckInst_3_n13 , \Check1_CheckInst_3_n12 ,
         \Check1_CheckInst_3_n11 , \Check1_CheckInst_3_n10 ,
         \Check1_CheckInst_3_n9 , \Check1_CheckInst_3_n8 ,
         \Check1_CheckInst_3_n7 , \Check1_CheckInst_3_n6 ,
         \Check1_CheckInst_3_n5 , \Check1_CheckInst_3_n4 ,
         \Check1_CheckInst_3_n3 ;
  wire   [63:0] MCOutput;
  wire   [63:0] AddRoundKeyOutput;
  wire   [63:0] PermutationOutput;
  wire   [63:0] Red_Input;
  wire   [63:0] Red_MCOutput;
  wire   [63:0] Red_K0;
  wire   [63:0] Red_AddRoundKeyOutput;
  wire   [63:0] Red_StateRegOutput;
  wire   [63:0] Red_Feedback;
  wire   [191:0] Red_SignaltoCheck;
  wire   [3:0] Error;

  NAND2_X1 \Check1_CheckInst_U9 ( .A1(Error[2]), .A2(Error[3]), .ZN(n9) );
  NAND2_X1 \Check1_CheckInst_U10 ( .A1(Error[0]), .A2(Error[1]), .ZN(n8) );
  OR2_X1 \Check1_CheckInst_U11 ( .A1(n9), .A2(n8), .ZN(ErrorFlag) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_0_U2  ( .A(\MCInst_XOR_r0_Inst_0_n3 ), .B(
        Input[0]), .ZN(MCOutput[48]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_0_U1  ( .A(Input[48]), .B(Input[16]), .ZN(
        \MCInst_XOR_r0_Inst_0_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_0_U1  ( .A(Input[32]), .B(Input[0]), .Z(
        MCOutput[32]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_1_U2  ( .A(\MCInst_XOR_r0_Inst_1_n3 ), .B(
        Input[1]), .ZN(MCOutput[49]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_1_U1  ( .A(Input[49]), .B(Input[17]), .ZN(
        \MCInst_XOR_r0_Inst_1_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_1_U1  ( .A(Input[33]), .B(Input[1]), .Z(
        MCOutput[33]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_2_U2  ( .A(\MCInst_XOR_r0_Inst_2_n3 ), .B(
        Input[2]), .ZN(MCOutput[50]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_2_U1  ( .A(Input[50]), .B(Input[18]), .ZN(
        \MCInst_XOR_r0_Inst_2_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_2_U1  ( .A(Input[34]), .B(Input[2]), .Z(
        MCOutput[34]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_3_U2  ( .A(\MCInst_XOR_r0_Inst_3_n3 ), .B(
        Input[3]), .ZN(MCOutput[51]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_3_U1  ( .A(Input[51]), .B(Input[19]), .ZN(
        \MCInst_XOR_r0_Inst_3_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_3_U1  ( .A(Input[35]), .B(Input[3]), .Z(
        MCOutput[35]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_4_U2  ( .A(\MCInst_XOR_r0_Inst_4_n3 ), .B(
        Input[4]), .ZN(MCOutput[52]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_4_U1  ( .A(Input[52]), .B(Input[20]), .ZN(
        \MCInst_XOR_r0_Inst_4_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_4_U1  ( .A(Input[36]), .B(Input[4]), .Z(
        MCOutput[36]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_5_U2  ( .A(\MCInst_XOR_r0_Inst_5_n3 ), .B(
        Input[5]), .ZN(MCOutput[53]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_5_U1  ( .A(Input[53]), .B(Input[21]), .ZN(
        \MCInst_XOR_r0_Inst_5_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_5_U1  ( .A(Input[37]), .B(Input[5]), .Z(
        MCOutput[37]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_6_U2  ( .A(\MCInst_XOR_r0_Inst_6_n3 ), .B(
        Input[6]), .ZN(MCOutput[54]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_6_U1  ( .A(Input[54]), .B(Input[22]), .ZN(
        \MCInst_XOR_r0_Inst_6_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_6_U1  ( .A(Input[38]), .B(Input[6]), .Z(
        MCOutput[38]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_7_U2  ( .A(\MCInst_XOR_r0_Inst_7_n3 ), .B(
        Input[7]), .ZN(MCOutput[55]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_7_U1  ( .A(Input[55]), .B(Input[23]), .ZN(
        \MCInst_XOR_r0_Inst_7_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_7_U1  ( .A(Input[39]), .B(Input[7]), .Z(
        MCOutput[39]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_8_U2  ( .A(\MCInst_XOR_r0_Inst_8_n3 ), .B(
        Input[8]), .ZN(MCOutput[56]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_8_U1  ( .A(Input[56]), .B(Input[24]), .ZN(
        \MCInst_XOR_r0_Inst_8_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_8_U1  ( .A(Input[40]), .B(Input[8]), .Z(
        MCOutput[40]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_9_U2  ( .A(\MCInst_XOR_r0_Inst_9_n3 ), .B(
        Input[9]), .ZN(MCOutput[57]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_9_U1  ( .A(Input[57]), .B(Input[25]), .ZN(
        \MCInst_XOR_r0_Inst_9_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_9_U1  ( .A(Input[41]), .B(Input[9]), .Z(
        MCOutput[41]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_10_U2  ( .A(\MCInst_XOR_r0_Inst_10_n3 ), .B(
        Input[10]), .ZN(MCOutput[58]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_10_U1  ( .A(Input[58]), .B(Input[26]), .ZN(
        \MCInst_XOR_r0_Inst_10_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_10_U1  ( .A(Input[42]), .B(Input[10]), .Z(
        MCOutput[42]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_11_U2  ( .A(\MCInst_XOR_r0_Inst_11_n3 ), .B(
        Input[11]), .ZN(MCOutput[59]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_11_U1  ( .A(Input[59]), .B(Input[27]), .ZN(
        \MCInst_XOR_r0_Inst_11_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_11_U1  ( .A(Input[43]), .B(Input[11]), .Z(
        MCOutput[43]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_12_U2  ( .A(\MCInst_XOR_r0_Inst_12_n3 ), .B(
        Input[12]), .ZN(MCOutput[60]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_12_U1  ( .A(Input[60]), .B(Input[28]), .ZN(
        \MCInst_XOR_r0_Inst_12_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_12_U1  ( .A(Input[44]), .B(Input[12]), .Z(
        MCOutput[44]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_13_U2  ( .A(\MCInst_XOR_r0_Inst_13_n3 ), .B(
        Input[13]), .ZN(MCOutput[61]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_13_U1  ( .A(Input[61]), .B(Input[29]), .ZN(
        \MCInst_XOR_r0_Inst_13_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_13_U1  ( .A(Input[45]), .B(Input[13]), .Z(
        MCOutput[45]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_14_U2  ( .A(\MCInst_XOR_r0_Inst_14_n3 ), .B(
        Input[14]), .ZN(MCOutput[62]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_14_U1  ( .A(Input[62]), .B(Input[30]), .ZN(
        \MCInst_XOR_r0_Inst_14_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_14_U1  ( .A(Input[46]), .B(Input[14]), .Z(
        MCOutput[46]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_15_U2  ( .A(\MCInst_XOR_r0_Inst_15_n3 ), .B(
        Input[15]), .ZN(MCOutput[63]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_15_U1  ( .A(Input[63]), .B(Input[31]), .ZN(
        \MCInst_XOR_r0_Inst_15_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_15_U1  ( .A(Input[47]), .B(Input[15]), .Z(
        MCOutput[47]) );
  XOR2_X1 \AddKeyXOR1_XORInst_0_0_U1  ( .A(MCOutput[48]), .B(Key[48]), .Z(
        AddRoundKeyOutput[48]) );
  XOR2_X1 \AddKeyXOR1_XORInst_0_1_U1  ( .A(MCOutput[49]), .B(Key[49]), .Z(
        AddRoundKeyOutput[49]) );
  XOR2_X1 \AddKeyXOR1_XORInst_0_2_U1  ( .A(MCOutput[50]), .B(Key[50]), .Z(
        AddRoundKeyOutput[50]) );
  XOR2_X1 \AddKeyXOR1_XORInst_0_3_U1  ( .A(MCOutput[51]), .B(Key[51]), .Z(
        AddRoundKeyOutput[51]) );
  XOR2_X1 \AddKeyXOR1_XORInst_1_0_U1  ( .A(MCOutput[52]), .B(Key[52]), .Z(
        AddRoundKeyOutput[52]) );
  XOR2_X1 \AddKeyXOR1_XORInst_1_1_U1  ( .A(MCOutput[53]), .B(Key[53]), .Z(
        AddRoundKeyOutput[53]) );
  XOR2_X1 \AddKeyXOR1_XORInst_1_2_U1  ( .A(MCOutput[54]), .B(Key[54]), .Z(
        AddRoundKeyOutput[54]) );
  XOR2_X1 \AddKeyXOR1_XORInst_1_3_U1  ( .A(MCOutput[55]), .B(Key[55]), .Z(
        AddRoundKeyOutput[55]) );
  XOR2_X1 \AddKeyXOR1_XORInst_2_0_U1  ( .A(MCOutput[56]), .B(Key[56]), .Z(
        AddRoundKeyOutput[56]) );
  XOR2_X1 \AddKeyXOR1_XORInst_2_1_U1  ( .A(MCOutput[57]), .B(Key[57]), .Z(
        AddRoundKeyOutput[57]) );
  XOR2_X1 \AddKeyXOR1_XORInst_2_2_U1  ( .A(MCOutput[58]), .B(Key[58]), .Z(
        AddRoundKeyOutput[58]) );
  XOR2_X1 \AddKeyXOR1_XORInst_2_3_U1  ( .A(MCOutput[59]), .B(Key[59]), .Z(
        AddRoundKeyOutput[59]) );
  XOR2_X1 \AddKeyXOR1_XORInst_3_0_U1  ( .A(MCOutput[60]), .B(Key[60]), .Z(
        AddRoundKeyOutput[60]) );
  XOR2_X1 \AddKeyXOR1_XORInst_3_1_U1  ( .A(MCOutput[61]), .B(Key[61]), .Z(
        AddRoundKeyOutput[61]) );
  XOR2_X1 \AddKeyXOR1_XORInst_3_2_U1  ( .A(MCOutput[62]), .B(Key[62]), .Z(
        AddRoundKeyOutput[62]) );
  XOR2_X1 \AddKeyXOR1_XORInst_3_3_U1  ( .A(MCOutput[63]), .B(Key[63]), .Z(
        AddRoundKeyOutput[63]) );
  XOR2_X1 \AddKeyConstXOR_XORInst_0_0_U1  ( .A(Key[40]), .B(MCOutput[40]), .Z(
        AddRoundKeyOutput[40]) );
  XOR2_X1 \AddKeyConstXOR_XORInst_0_1_U1  ( .A(Key[41]), .B(MCOutput[41]), .Z(
        AddRoundKeyOutput[41]) );
  XOR2_X1 \AddKeyConstXOR_XORInst_0_2_U1  ( .A(Key[42]), .B(MCOutput[42]), .Z(
        AddRoundKeyOutput[42]) );
  XOR2_X1 \AddKeyConstXOR_XORInst_0_3_U1  ( .A(Key[43]), .B(MCOutput[43]), .Z(
        AddRoundKeyOutput[43]) );
  XOR2_X1 \AddKeyConstXOR_XORInst_1_0_U1  ( .A(Key[44]), .B(MCOutput[44]), .Z(
        AddRoundKeyOutput[44]) );
  XOR2_X1 \AddKeyConstXOR_XORInst_1_1_U1  ( .A(Key[45]), .B(MCOutput[45]), .Z(
        AddRoundKeyOutput[45]) );
  XOR2_X1 \AddKeyConstXOR_XORInst_1_2_U1  ( .A(Key[46]), .B(MCOutput[46]), .Z(
        AddRoundKeyOutput[46]) );
  XOR2_X1 \AddKeyConstXOR_XORInst_1_3_U1  ( .A(Key[47]), .B(MCOutput[47]), .Z(
        AddRoundKeyOutput[47]) );
  XOR2_X1 \AddKeyXOR2_XORInst_0_0_U1  ( .A(Input[0]), .B(Key[0]), .Z(
        AddRoundKeyOutput[0]) );
  XOR2_X1 \AddKeyXOR2_XORInst_0_1_U1  ( .A(Input[1]), .B(Key[1]), .Z(
        AddRoundKeyOutput[1]) );
  XOR2_X1 \AddKeyXOR2_XORInst_0_2_U1  ( .A(Input[2]), .B(Key[2]), .Z(
        AddRoundKeyOutput[2]) );
  XOR2_X1 \AddKeyXOR2_XORInst_0_3_U1  ( .A(Input[3]), .B(Key[3]), .Z(
        AddRoundKeyOutput[3]) );
  XOR2_X1 \AddKeyXOR2_XORInst_1_0_U1  ( .A(Input[4]), .B(Key[4]), .Z(
        AddRoundKeyOutput[4]) );
  XOR2_X1 \AddKeyXOR2_XORInst_1_1_U1  ( .A(Input[5]), .B(Key[5]), .Z(
        AddRoundKeyOutput[5]) );
  XOR2_X1 \AddKeyXOR2_XORInst_1_2_U1  ( .A(Input[6]), .B(Key[6]), .Z(
        AddRoundKeyOutput[6]) );
  XOR2_X1 \AddKeyXOR2_XORInst_1_3_U1  ( .A(Input[7]), .B(Key[7]), .Z(
        AddRoundKeyOutput[7]) );
  XOR2_X1 \AddKeyXOR2_XORInst_2_0_U1  ( .A(Input[8]), .B(Key[8]), .Z(
        AddRoundKeyOutput[8]) );
  XOR2_X1 \AddKeyXOR2_XORInst_2_1_U1  ( .A(Input[9]), .B(Key[9]), .Z(
        AddRoundKeyOutput[9]) );
  XOR2_X1 \AddKeyXOR2_XORInst_2_2_U1  ( .A(Input[10]), .B(Key[10]), .Z(
        AddRoundKeyOutput[10]) );
  XOR2_X1 \AddKeyXOR2_XORInst_2_3_U1  ( .A(Input[11]), .B(Key[11]), .Z(
        AddRoundKeyOutput[11]) );
  XOR2_X1 \AddKeyXOR2_XORInst_3_0_U1  ( .A(Input[12]), .B(Key[12]), .Z(
        AddRoundKeyOutput[12]) );
  XOR2_X1 \AddKeyXOR2_XORInst_3_1_U1  ( .A(Input[13]), .B(Key[13]), .Z(
        AddRoundKeyOutput[13]) );
  XOR2_X1 \AddKeyXOR2_XORInst_3_2_U1  ( .A(Input[14]), .B(Key[14]), .Z(
        AddRoundKeyOutput[14]) );
  XOR2_X1 \AddKeyXOR2_XORInst_3_3_U1  ( .A(Input[15]), .B(Key[15]), .Z(
        AddRoundKeyOutput[15]) );
  XOR2_X1 \AddKeyXOR2_XORInst_4_0_U1  ( .A(Input[16]), .B(Key[16]), .Z(
        AddRoundKeyOutput[16]) );
  XOR2_X1 \AddKeyXOR2_XORInst_4_1_U1  ( .A(Input[17]), .B(Key[17]), .Z(
        AddRoundKeyOutput[17]) );
  XOR2_X1 \AddKeyXOR2_XORInst_4_2_U1  ( .A(Input[18]), .B(Key[18]), .Z(
        AddRoundKeyOutput[18]) );
  XOR2_X1 \AddKeyXOR2_XORInst_4_3_U1  ( .A(Input[19]), .B(Key[19]), .Z(
        AddRoundKeyOutput[19]) );
  XOR2_X1 \AddKeyXOR2_XORInst_5_0_U1  ( .A(Input[20]), .B(Key[20]), .Z(
        AddRoundKeyOutput[20]) );
  XOR2_X1 \AddKeyXOR2_XORInst_5_1_U1  ( .A(Input[21]), .B(Key[21]), .Z(
        AddRoundKeyOutput[21]) );
  XOR2_X1 \AddKeyXOR2_XORInst_5_2_U1  ( .A(Input[22]), .B(Key[22]), .Z(
        AddRoundKeyOutput[22]) );
  XOR2_X1 \AddKeyXOR2_XORInst_5_3_U1  ( .A(Input[23]), .B(Key[23]), .Z(
        AddRoundKeyOutput[23]) );
  XOR2_X1 \AddKeyXOR2_XORInst_6_0_U1  ( .A(Input[24]), .B(Key[24]), .Z(
        AddRoundKeyOutput[24]) );
  XOR2_X1 \AddKeyXOR2_XORInst_6_1_U1  ( .A(Input[25]), .B(Key[25]), .Z(
        AddRoundKeyOutput[25]) );
  XOR2_X1 \AddKeyXOR2_XORInst_6_2_U1  ( .A(Input[26]), .B(Key[26]), .Z(
        AddRoundKeyOutput[26]) );
  XOR2_X1 \AddKeyXOR2_XORInst_6_3_U1  ( .A(Input[27]), .B(Key[27]), .Z(
        AddRoundKeyOutput[27]) );
  XOR2_X1 \AddKeyXOR2_XORInst_7_0_U1  ( .A(Input[28]), .B(Key[28]), .Z(
        AddRoundKeyOutput[28]) );
  XOR2_X1 \AddKeyXOR2_XORInst_7_1_U1  ( .A(Input[29]), .B(Key[29]), .Z(
        AddRoundKeyOutput[29]) );
  XOR2_X1 \AddKeyXOR2_XORInst_7_2_U1  ( .A(Input[30]), .B(Key[30]), .Z(
        AddRoundKeyOutput[30]) );
  XOR2_X1 \AddKeyXOR2_XORInst_7_3_U1  ( .A(Input[31]), .B(Key[31]), .Z(
        AddRoundKeyOutput[31]) );
  XOR2_X1 \AddKeyXOR2_XORInst_8_0_U1  ( .A(MCOutput[32]), .B(Key[32]), .Z(
        AddRoundKeyOutput[32]) );
  XOR2_X1 \AddKeyXOR2_XORInst_8_1_U1  ( .A(MCOutput[33]), .B(Key[33]), .Z(
        AddRoundKeyOutput[33]) );
  XOR2_X1 \AddKeyXOR2_XORInst_8_2_U1  ( .A(MCOutput[34]), .B(Key[34]), .Z(
        AddRoundKeyOutput[34]) );
  XOR2_X1 \AddKeyXOR2_XORInst_8_3_U1  ( .A(MCOutput[35]), .B(Key[35]), .Z(
        AddRoundKeyOutput[35]) );
  XOR2_X1 \AddKeyXOR2_XORInst_9_0_U1  ( .A(MCOutput[36]), .B(Key[36]), .Z(
        AddRoundKeyOutput[36]) );
  XOR2_X1 \AddKeyXOR2_XORInst_9_1_U1  ( .A(MCOutput[37]), .B(Key[37]), .Z(
        AddRoundKeyOutput[37]) );
  XOR2_X1 \AddKeyXOR2_XORInst_9_2_U1  ( .A(MCOutput[38]), .B(Key[38]), .Z(
        AddRoundKeyOutput[38]) );
  XOR2_X1 \AddKeyXOR2_XORInst_9_3_U1  ( .A(MCOutput[39]), .B(Key[39]), .Z(
        AddRoundKeyOutput[39]) );
  DFF_X1 \StateReg_s_current_state_reg[0]  ( .D(AddRoundKeyOutput[0]), .CK(clk), .Q(PermutationOutput[60]) );
  DFF_X1 \StateReg_s_current_state_reg[1]  ( .D(AddRoundKeyOutput[1]), .CK(clk), .Q(PermutationOutput[61]) );
  DFF_X1 \StateReg_s_current_state_reg[2]  ( .D(AddRoundKeyOutput[2]), .CK(clk), .Q(PermutationOutput[62]) );
  DFF_X1 \StateReg_s_current_state_reg[3]  ( .D(AddRoundKeyOutput[3]), .CK(clk), .Q(PermutationOutput[63]) );
  DFF_X1 \StateReg_s_current_state_reg[4]  ( .D(AddRoundKeyOutput[4]), .CK(clk), .Q(PermutationOutput[48]) );
  DFF_X1 \StateReg_s_current_state_reg[5]  ( .D(AddRoundKeyOutput[5]), .CK(clk), .Q(PermutationOutput[49]) );
  DFF_X1 \StateReg_s_current_state_reg[6]  ( .D(AddRoundKeyOutput[6]), .CK(clk), .Q(PermutationOutput[50]) );
  DFF_X1 \StateReg_s_current_state_reg[7]  ( .D(AddRoundKeyOutput[7]), .CK(clk), .Q(PermutationOutput[51]) );
  DFF_X1 \StateReg_s_current_state_reg[8]  ( .D(AddRoundKeyOutput[8]), .CK(clk), .Q(PermutationOutput[52]) );
  DFF_X1 \StateReg_s_current_state_reg[9]  ( .D(AddRoundKeyOutput[9]), .CK(clk), .Q(PermutationOutput[53]) );
  DFF_X1 \StateReg_s_current_state_reg[10]  ( .D(AddRoundKeyOutput[10]), .CK(
        clk), .Q(PermutationOutput[54]) );
  DFF_X1 \StateReg_s_current_state_reg[11]  ( .D(AddRoundKeyOutput[11]), .CK(
        clk), .Q(PermutationOutput[55]) );
  DFF_X1 \StateReg_s_current_state_reg[12]  ( .D(AddRoundKeyOutput[12]), .CK(
        clk), .Q(PermutationOutput[56]) );
  DFF_X1 \StateReg_s_current_state_reg[13]  ( .D(AddRoundKeyOutput[13]), .CK(
        clk), .Q(PermutationOutput[57]) );
  DFF_X1 \StateReg_s_current_state_reg[14]  ( .D(AddRoundKeyOutput[14]), .CK(
        clk), .Q(PermutationOutput[58]) );
  DFF_X1 \StateReg_s_current_state_reg[15]  ( .D(AddRoundKeyOutput[15]), .CK(
        clk), .Q(PermutationOutput[59]) );
  DFF_X1 \StateReg_s_current_state_reg[16]  ( .D(AddRoundKeyOutput[16]), .CK(
        clk), .Q(PermutationOutput[32]) );
  DFF_X1 \StateReg_s_current_state_reg[17]  ( .D(AddRoundKeyOutput[17]), .CK(
        clk), .Q(PermutationOutput[33]) );
  DFF_X1 \StateReg_s_current_state_reg[18]  ( .D(AddRoundKeyOutput[18]), .CK(
        clk), .Q(PermutationOutput[34]) );
  DFF_X1 \StateReg_s_current_state_reg[19]  ( .D(AddRoundKeyOutput[19]), .CK(
        clk), .Q(PermutationOutput[35]) );
  DFF_X1 \StateReg_s_current_state_reg[20]  ( .D(AddRoundKeyOutput[20]), .CK(
        clk), .Q(PermutationOutput[44]) );
  DFF_X1 \StateReg_s_current_state_reg[21]  ( .D(AddRoundKeyOutput[21]), .CK(
        clk), .Q(PermutationOutput[45]) );
  DFF_X1 \StateReg_s_current_state_reg[22]  ( .D(AddRoundKeyOutput[22]), .CK(
        clk), .Q(PermutationOutput[46]) );
  DFF_X1 \StateReg_s_current_state_reg[23]  ( .D(AddRoundKeyOutput[23]), .CK(
        clk), .Q(PermutationOutput[47]) );
  DFF_X1 \StateReg_s_current_state_reg[24]  ( .D(AddRoundKeyOutput[24]), .CK(
        clk), .Q(PermutationOutput[40]) );
  DFF_X1 \StateReg_s_current_state_reg[25]  ( .D(AddRoundKeyOutput[25]), .CK(
        clk), .Q(PermutationOutput[41]) );
  DFF_X1 \StateReg_s_current_state_reg[26]  ( .D(AddRoundKeyOutput[26]), .CK(
        clk), .Q(PermutationOutput[42]) );
  DFF_X1 \StateReg_s_current_state_reg[27]  ( .D(AddRoundKeyOutput[27]), .CK(
        clk), .Q(PermutationOutput[43]) );
  DFF_X1 \StateReg_s_current_state_reg[28]  ( .D(AddRoundKeyOutput[28]), .CK(
        clk), .Q(PermutationOutput[36]) );
  DFF_X1 \StateReg_s_current_state_reg[29]  ( .D(AddRoundKeyOutput[29]), .CK(
        clk), .Q(PermutationOutput[37]) );
  DFF_X1 \StateReg_s_current_state_reg[30]  ( .D(AddRoundKeyOutput[30]), .CK(
        clk), .Q(PermutationOutput[38]) );
  DFF_X1 \StateReg_s_current_state_reg[31]  ( .D(AddRoundKeyOutput[31]), .CK(
        clk), .Q(PermutationOutput[39]) );
  DFF_X1 \StateReg_s_current_state_reg[32]  ( .D(AddRoundKeyOutput[32]), .CK(
        clk), .Q(PermutationOutput[16]) );
  DFF_X1 \StateReg_s_current_state_reg[33]  ( .D(AddRoundKeyOutput[33]), .CK(
        clk), .Q(PermutationOutput[17]) );
  DFF_X1 \StateReg_s_current_state_reg[34]  ( .D(AddRoundKeyOutput[34]), .CK(
        clk), .Q(PermutationOutput[18]) );
  DFF_X1 \StateReg_s_current_state_reg[35]  ( .D(AddRoundKeyOutput[35]), .CK(
        clk), .Q(PermutationOutput[19]) );
  DFF_X1 \StateReg_s_current_state_reg[36]  ( .D(AddRoundKeyOutput[36]), .CK(
        clk), .Q(PermutationOutput[28]) );
  DFF_X1 \StateReg_s_current_state_reg[37]  ( .D(AddRoundKeyOutput[37]), .CK(
        clk), .Q(PermutationOutput[29]) );
  DFF_X1 \StateReg_s_current_state_reg[38]  ( .D(AddRoundKeyOutput[38]), .CK(
        clk), .Q(PermutationOutput[30]) );
  DFF_X1 \StateReg_s_current_state_reg[39]  ( .D(AddRoundKeyOutput[39]), .CK(
        clk), .Q(PermutationOutput[31]) );
  DFF_X1 \StateReg_s_current_state_reg[40]  ( .D(AddRoundKeyOutput[40]), .CK(
        clk), .Q(PermutationOutput[24]) );
  DFF_X1 \StateReg_s_current_state_reg[41]  ( .D(AddRoundKeyOutput[41]), .CK(
        clk), .Q(PermutationOutput[25]) );
  DFF_X1 \StateReg_s_current_state_reg[42]  ( .D(AddRoundKeyOutput[42]), .CK(
        clk), .Q(PermutationOutput[26]) );
  DFF_X1 \StateReg_s_current_state_reg[43]  ( .D(AddRoundKeyOutput[43]), .CK(
        clk), .Q(PermutationOutput[27]) );
  DFF_X1 \StateReg_s_current_state_reg[44]  ( .D(AddRoundKeyOutput[44]), .CK(
        clk), .Q(PermutationOutput[20]) );
  DFF_X1 \StateReg_s_current_state_reg[45]  ( .D(AddRoundKeyOutput[45]), .CK(
        clk), .Q(PermutationOutput[21]) );
  DFF_X1 \StateReg_s_current_state_reg[46]  ( .D(AddRoundKeyOutput[46]), .CK(
        clk), .Q(PermutationOutput[22]) );
  DFF_X1 \StateReg_s_current_state_reg[47]  ( .D(AddRoundKeyOutput[47]), .CK(
        clk), .Q(PermutationOutput[23]) );
  DFF_X1 \StateReg_s_current_state_reg[48]  ( .D(AddRoundKeyOutput[48]), .CK(
        clk), .Q(PermutationOutput[4]) );
  DFF_X1 \StateReg_s_current_state_reg[49]  ( .D(AddRoundKeyOutput[49]), .CK(
        clk), .Q(PermutationOutput[5]) );
  DFF_X1 \StateReg_s_current_state_reg[50]  ( .D(AddRoundKeyOutput[50]), .CK(
        clk), .Q(PermutationOutput[6]) );
  DFF_X1 \StateReg_s_current_state_reg[51]  ( .D(AddRoundKeyOutput[51]), .CK(
        clk), .Q(PermutationOutput[7]) );
  DFF_X1 \StateReg_s_current_state_reg[52]  ( .D(AddRoundKeyOutput[52]), .CK(
        clk), .Q(PermutationOutput[8]) );
  DFF_X1 \StateReg_s_current_state_reg[53]  ( .D(AddRoundKeyOutput[53]), .CK(
        clk), .Q(PermutationOutput[9]) );
  DFF_X1 \StateReg_s_current_state_reg[54]  ( .D(AddRoundKeyOutput[54]), .CK(
        clk), .Q(PermutationOutput[10]) );
  DFF_X1 \StateReg_s_current_state_reg[55]  ( .D(AddRoundKeyOutput[55]), .CK(
        clk), .Q(PermutationOutput[11]) );
  DFF_X1 \StateReg_s_current_state_reg[56]  ( .D(AddRoundKeyOutput[56]), .CK(
        clk), .Q(PermutationOutput[12]) );
  DFF_X1 \StateReg_s_current_state_reg[57]  ( .D(AddRoundKeyOutput[57]), .CK(
        clk), .Q(PermutationOutput[13]) );
  DFF_X1 \StateReg_s_current_state_reg[58]  ( .D(AddRoundKeyOutput[58]), .CK(
        clk), .Q(PermutationOutput[14]) );
  DFF_X1 \StateReg_s_current_state_reg[59]  ( .D(AddRoundKeyOutput[59]), .CK(
        clk), .Q(PermutationOutput[15]) );
  DFF_X1 \StateReg_s_current_state_reg[60]  ( .D(AddRoundKeyOutput[60]), .CK(
        clk), .Q(PermutationOutput[0]) );
  DFF_X1 \StateReg_s_current_state_reg[61]  ( .D(AddRoundKeyOutput[61]), .CK(
        clk), .Q(PermutationOutput[1]) );
  DFF_X1 \StateReg_s_current_state_reg[62]  ( .D(AddRoundKeyOutput[62]), .CK(
        clk), .Q(PermutationOutput[2]) );
  DFF_X1 \StateReg_s_current_state_reg[63]  ( .D(AddRoundKeyOutput[63]), .CK(
        clk), .Q(PermutationOutput[3]) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_0_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_0_LFInst_0_n10 ), .ZN(Output[0]) );
  AND2_X1 \SubCellInst_LFInst_0_LFInst_0_U7  ( .A1(PermutationOutput[3]), .A2(
        PermutationOutput[2]), .ZN(\SubCellInst_LFInst_0_LFInst_0_n10 ) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_0_U6  ( .A1(PermutationOutput[1]), .A2(
        \SubCellInst_LFInst_0_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_0_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_0_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_0_U4  ( .A1(PermutationOutput[3]), .A2(
        PermutationOutput[2]), .ZN(\SubCellInst_LFInst_0_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_0_LFInst_0_U3  ( .A(PermutationOutput[0]), .ZN(
        \SubCellInst_LFInst_0_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_0_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_0_LFInst_1_n5 ), .ZN(Output[1]) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U5  ( .A1(PermutationOutput[2]), 
        .A2(PermutationOutput[0]), .ZN(\SubCellInst_LFInst_0_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_0_LFInst_1_U4  ( .A1(PermutationOutput[3]), .A2(
        \SubCellInst_LFInst_0_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_1_U3  ( .A1(PermutationOutput[2]), .A2(
        PermutationOutput[0]), .ZN(\SubCellInst_LFInst_0_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_0_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_0_LFInst_2_n10 ), .ZN(Output[2]) );
  OR2_X1 \SubCellInst_LFInst_0_LFInst_2_U7  ( .A1(PermutationOutput[0]), .A2(
        PermutationOutput[3]), .ZN(\SubCellInst_LFInst_0_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U6  ( .A1(PermutationOutput[1]), 
        .A2(\SubCellInst_LFInst_0_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_0_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_0_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U4  ( .A1(PermutationOutput[0]), 
        .A2(PermutationOutput[3]), .ZN(\SubCellInst_LFInst_0_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_0_LFInst_2_U3  ( .A(PermutationOutput[2]), .ZN(
        \SubCellInst_LFInst_0_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_0_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_0_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_0_LFInst_3_n5 ), .ZN(Output[3]) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_3_U5  ( .A1(PermutationOutput[3]), .A2(
        PermutationOutput[0]), .ZN(\SubCellInst_LFInst_0_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_3_U4  ( .A1(PermutationOutput[1]), .A2(
        \SubCellInst_LFInst_0_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_0_LFInst_3_U3  ( .A1(PermutationOutput[3]), .A2(
        PermutationOutput[2]), .ZN(\SubCellInst_LFInst_0_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_1_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_1_LFInst_0_n10 ), .ZN(Output[4]) );
  AND2_X1 \SubCellInst_LFInst_1_LFInst_0_U7  ( .A1(PermutationOutput[7]), .A2(
        PermutationOutput[6]), .ZN(\SubCellInst_LFInst_1_LFInst_0_n10 ) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_0_U6  ( .A1(PermutationOutput[5]), .A2(
        \SubCellInst_LFInst_1_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_1_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_1_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_0_U4  ( .A1(PermutationOutput[7]), .A2(
        PermutationOutput[6]), .ZN(\SubCellInst_LFInst_1_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_1_LFInst_0_U3  ( .A(PermutationOutput[4]), .ZN(
        \SubCellInst_LFInst_1_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_1_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_1_LFInst_1_n5 ), .ZN(Output[5]) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U5  ( .A1(PermutationOutput[6]), 
        .A2(PermutationOutput[4]), .ZN(\SubCellInst_LFInst_1_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_1_LFInst_1_U4  ( .A1(PermutationOutput[7]), .A2(
        \SubCellInst_LFInst_1_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_1_U3  ( .A1(PermutationOutput[6]), .A2(
        PermutationOutput[4]), .ZN(\SubCellInst_LFInst_1_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_1_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_1_LFInst_2_n10 ), .ZN(Output[6]) );
  OR2_X1 \SubCellInst_LFInst_1_LFInst_2_U7  ( .A1(PermutationOutput[4]), .A2(
        PermutationOutput[7]), .ZN(\SubCellInst_LFInst_1_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U6  ( .A1(PermutationOutput[5]), 
        .A2(\SubCellInst_LFInst_1_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_1_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_1_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U4  ( .A1(PermutationOutput[4]), 
        .A2(PermutationOutput[7]), .ZN(\SubCellInst_LFInst_1_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_1_LFInst_2_U3  ( .A(PermutationOutput[6]), .ZN(
        \SubCellInst_LFInst_1_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_1_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_1_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_1_LFInst_3_n5 ), .ZN(Output[7]) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_3_U5  ( .A1(PermutationOutput[7]), .A2(
        PermutationOutput[4]), .ZN(\SubCellInst_LFInst_1_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_3_U4  ( .A1(PermutationOutput[5]), .A2(
        \SubCellInst_LFInst_1_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_1_LFInst_3_U3  ( .A1(PermutationOutput[7]), .A2(
        PermutationOutput[6]), .ZN(\SubCellInst_LFInst_1_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_2_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_2_LFInst_0_n10 ), .ZN(Output[8]) );
  AND2_X1 \SubCellInst_LFInst_2_LFInst_0_U7  ( .A1(PermutationOutput[11]), 
        .A2(PermutationOutput[10]), .ZN(\SubCellInst_LFInst_2_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_0_U6  ( .A1(PermutationOutput[9]), .A2(
        \SubCellInst_LFInst_2_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_2_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_2_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_0_U4  ( .A1(PermutationOutput[11]), 
        .A2(PermutationOutput[10]), .ZN(\SubCellInst_LFInst_2_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_2_LFInst_0_U3  ( .A(PermutationOutput[8]), .ZN(
        \SubCellInst_LFInst_2_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_2_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_2_LFInst_1_n5 ), .ZN(Output[9]) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U5  ( .A1(PermutationOutput[10]), 
        .A2(PermutationOutput[8]), .ZN(\SubCellInst_LFInst_2_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_2_LFInst_1_U4  ( .A1(PermutationOutput[11]), .A2(
        \SubCellInst_LFInst_2_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_1_U3  ( .A1(PermutationOutput[10]), 
        .A2(PermutationOutput[8]), .ZN(\SubCellInst_LFInst_2_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_2_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_2_LFInst_2_n10 ), .ZN(Output[10]) );
  OR2_X1 \SubCellInst_LFInst_2_LFInst_2_U7  ( .A1(PermutationOutput[8]), .A2(
        PermutationOutput[11]), .ZN(\SubCellInst_LFInst_2_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U6  ( .A1(PermutationOutput[9]), 
        .A2(\SubCellInst_LFInst_2_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_2_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_2_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U4  ( .A1(PermutationOutput[8]), 
        .A2(PermutationOutput[11]), .ZN(\SubCellInst_LFInst_2_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_2_LFInst_2_U3  ( .A(PermutationOutput[10]), .ZN(
        \SubCellInst_LFInst_2_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_2_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_2_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_2_LFInst_3_n5 ), .ZN(Output[11]) );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_3_U5  ( .A1(PermutationOutput[11]), 
        .A2(PermutationOutput[8]), .ZN(\SubCellInst_LFInst_2_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_3_U4  ( .A1(PermutationOutput[9]), .A2(
        \SubCellInst_LFInst_2_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_2_LFInst_3_U3  ( .A1(PermutationOutput[11]), 
        .A2(PermutationOutput[10]), .ZN(\SubCellInst_LFInst_2_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_3_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_3_LFInst_0_n10 ), .ZN(Output[12]) );
  AND2_X1 \SubCellInst_LFInst_3_LFInst_0_U7  ( .A1(PermutationOutput[15]), 
        .A2(PermutationOutput[14]), .ZN(\SubCellInst_LFInst_3_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_0_U6  ( .A1(PermutationOutput[13]), 
        .A2(\SubCellInst_LFInst_3_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_3_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_3_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_0_U4  ( .A1(PermutationOutput[15]), 
        .A2(PermutationOutput[14]), .ZN(\SubCellInst_LFInst_3_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_3_LFInst_0_U3  ( .A(PermutationOutput[12]), .ZN(
        \SubCellInst_LFInst_3_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_3_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_3_LFInst_1_n5 ), .ZN(Output[13]) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U5  ( .A1(PermutationOutput[14]), 
        .A2(PermutationOutput[12]), .ZN(\SubCellInst_LFInst_3_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_3_LFInst_1_U4  ( .A1(PermutationOutput[15]), .A2(
        \SubCellInst_LFInst_3_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_1_U3  ( .A1(PermutationOutput[14]), 
        .A2(PermutationOutput[12]), .ZN(\SubCellInst_LFInst_3_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_3_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_3_LFInst_2_n10 ), .ZN(Output[14]) );
  OR2_X1 \SubCellInst_LFInst_3_LFInst_2_U7  ( .A1(PermutationOutput[12]), .A2(
        PermutationOutput[15]), .ZN(\SubCellInst_LFInst_3_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U6  ( .A1(PermutationOutput[13]), 
        .A2(\SubCellInst_LFInst_3_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_3_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_3_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U4  ( .A1(PermutationOutput[12]), 
        .A2(PermutationOutput[15]), .ZN(\SubCellInst_LFInst_3_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_3_LFInst_2_U3  ( .A(PermutationOutput[14]), .ZN(
        \SubCellInst_LFInst_3_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_3_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_3_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_3_LFInst_3_n5 ), .ZN(Output[15]) );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_3_U5  ( .A1(PermutationOutput[15]), 
        .A2(PermutationOutput[12]), .ZN(\SubCellInst_LFInst_3_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_3_U4  ( .A1(PermutationOutput[13]), 
        .A2(\SubCellInst_LFInst_3_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_3_LFInst_3_U3  ( .A1(PermutationOutput[15]), 
        .A2(PermutationOutput[14]), .ZN(\SubCellInst_LFInst_3_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_4_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_4_LFInst_0_n10 ), .ZN(Output[16]) );
  AND2_X1 \SubCellInst_LFInst_4_LFInst_0_U7  ( .A1(PermutationOutput[19]), 
        .A2(PermutationOutput[18]), .ZN(\SubCellInst_LFInst_4_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_0_U6  ( .A1(PermutationOutput[17]), 
        .A2(\SubCellInst_LFInst_4_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_4_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_4_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_0_U4  ( .A1(PermutationOutput[19]), 
        .A2(PermutationOutput[18]), .ZN(\SubCellInst_LFInst_4_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_4_LFInst_0_U3  ( .A(PermutationOutput[16]), .ZN(
        \SubCellInst_LFInst_4_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_4_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_4_LFInst_1_n5 ), .ZN(Output[17]) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U5  ( .A1(PermutationOutput[18]), 
        .A2(PermutationOutput[16]), .ZN(\SubCellInst_LFInst_4_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_4_LFInst_1_U4  ( .A1(PermutationOutput[19]), .A2(
        \SubCellInst_LFInst_4_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_1_U3  ( .A1(PermutationOutput[18]), 
        .A2(PermutationOutput[16]), .ZN(\SubCellInst_LFInst_4_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_4_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_4_LFInst_2_n10 ), .ZN(Output[18]) );
  OR2_X1 \SubCellInst_LFInst_4_LFInst_2_U7  ( .A1(PermutationOutput[16]), .A2(
        PermutationOutput[19]), .ZN(\SubCellInst_LFInst_4_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U6  ( .A1(PermutationOutput[17]), 
        .A2(\SubCellInst_LFInst_4_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_4_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_4_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U4  ( .A1(PermutationOutput[16]), 
        .A2(PermutationOutput[19]), .ZN(\SubCellInst_LFInst_4_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_4_LFInst_2_U3  ( .A(PermutationOutput[18]), .ZN(
        \SubCellInst_LFInst_4_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_4_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_4_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_4_LFInst_3_n5 ), .ZN(Output[19]) );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_3_U5  ( .A1(PermutationOutput[19]), 
        .A2(PermutationOutput[16]), .ZN(\SubCellInst_LFInst_4_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_3_U4  ( .A1(PermutationOutput[17]), 
        .A2(\SubCellInst_LFInst_4_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_4_LFInst_3_U3  ( .A1(PermutationOutput[19]), 
        .A2(PermutationOutput[18]), .ZN(\SubCellInst_LFInst_4_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_5_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_5_LFInst_0_n10 ), .ZN(Output[20]) );
  AND2_X1 \SubCellInst_LFInst_5_LFInst_0_U7  ( .A1(PermutationOutput[23]), 
        .A2(PermutationOutput[22]), .ZN(\SubCellInst_LFInst_5_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_0_U6  ( .A1(PermutationOutput[21]), 
        .A2(\SubCellInst_LFInst_5_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_5_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_5_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_0_U4  ( .A1(PermutationOutput[23]), 
        .A2(PermutationOutput[22]), .ZN(\SubCellInst_LFInst_5_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_5_LFInst_0_U3  ( .A(PermutationOutput[20]), .ZN(
        \SubCellInst_LFInst_5_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_5_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_5_LFInst_1_n5 ), .ZN(Output[21]) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U5  ( .A1(PermutationOutput[22]), 
        .A2(PermutationOutput[20]), .ZN(\SubCellInst_LFInst_5_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_5_LFInst_1_U4  ( .A1(PermutationOutput[23]), .A2(
        \SubCellInst_LFInst_5_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_1_U3  ( .A1(PermutationOutput[22]), 
        .A2(PermutationOutput[20]), .ZN(\SubCellInst_LFInst_5_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_5_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_5_LFInst_2_n10 ), .ZN(Output[22]) );
  OR2_X1 \SubCellInst_LFInst_5_LFInst_2_U7  ( .A1(PermutationOutput[20]), .A2(
        PermutationOutput[23]), .ZN(\SubCellInst_LFInst_5_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U6  ( .A1(PermutationOutput[21]), 
        .A2(\SubCellInst_LFInst_5_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_5_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_5_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U4  ( .A1(PermutationOutput[20]), 
        .A2(PermutationOutput[23]), .ZN(\SubCellInst_LFInst_5_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_5_LFInst_2_U3  ( .A(PermutationOutput[22]), .ZN(
        \SubCellInst_LFInst_5_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_5_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_5_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_5_LFInst_3_n5 ), .ZN(Output[23]) );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_3_U5  ( .A1(PermutationOutput[23]), 
        .A2(PermutationOutput[20]), .ZN(\SubCellInst_LFInst_5_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_3_U4  ( .A1(PermutationOutput[21]), 
        .A2(\SubCellInst_LFInst_5_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_5_LFInst_3_U3  ( .A1(PermutationOutput[23]), 
        .A2(PermutationOutput[22]), .ZN(\SubCellInst_LFInst_5_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_6_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_6_LFInst_0_n10 ), .ZN(Output[24]) );
  AND2_X1 \SubCellInst_LFInst_6_LFInst_0_U7  ( .A1(PermutationOutput[27]), 
        .A2(PermutationOutput[26]), .ZN(\SubCellInst_LFInst_6_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_0_U6  ( .A1(PermutationOutput[25]), 
        .A2(\SubCellInst_LFInst_6_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_6_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_6_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_0_U4  ( .A1(PermutationOutput[27]), 
        .A2(PermutationOutput[26]), .ZN(\SubCellInst_LFInst_6_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_6_LFInst_0_U3  ( .A(PermutationOutput[24]), .ZN(
        \SubCellInst_LFInst_6_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_6_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_6_LFInst_1_n5 ), .ZN(Output[25]) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U5  ( .A1(PermutationOutput[26]), 
        .A2(PermutationOutput[24]), .ZN(\SubCellInst_LFInst_6_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_6_LFInst_1_U4  ( .A1(PermutationOutput[27]), .A2(
        \SubCellInst_LFInst_6_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_1_U3  ( .A1(PermutationOutput[26]), 
        .A2(PermutationOutput[24]), .ZN(\SubCellInst_LFInst_6_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_6_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_6_LFInst_2_n10 ), .ZN(Output[26]) );
  OR2_X1 \SubCellInst_LFInst_6_LFInst_2_U7  ( .A1(PermutationOutput[24]), .A2(
        PermutationOutput[27]), .ZN(\SubCellInst_LFInst_6_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U6  ( .A1(PermutationOutput[25]), 
        .A2(\SubCellInst_LFInst_6_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_6_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_6_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U4  ( .A1(PermutationOutput[24]), 
        .A2(PermutationOutput[27]), .ZN(\SubCellInst_LFInst_6_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_6_LFInst_2_U3  ( .A(PermutationOutput[26]), .ZN(
        \SubCellInst_LFInst_6_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_6_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_6_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_6_LFInst_3_n5 ), .ZN(Output[27]) );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_3_U5  ( .A1(PermutationOutput[27]), 
        .A2(PermutationOutput[24]), .ZN(\SubCellInst_LFInst_6_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_3_U4  ( .A1(PermutationOutput[25]), 
        .A2(\SubCellInst_LFInst_6_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_6_LFInst_3_U3  ( .A1(PermutationOutput[27]), 
        .A2(PermutationOutput[26]), .ZN(\SubCellInst_LFInst_6_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_7_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_7_LFInst_0_n10 ), .ZN(Output[28]) );
  AND2_X1 \SubCellInst_LFInst_7_LFInst_0_U7  ( .A1(PermutationOutput[31]), 
        .A2(PermutationOutput[30]), .ZN(\SubCellInst_LFInst_7_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_0_U6  ( .A1(PermutationOutput[29]), 
        .A2(\SubCellInst_LFInst_7_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_7_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_7_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_0_U4  ( .A1(PermutationOutput[31]), 
        .A2(PermutationOutput[30]), .ZN(\SubCellInst_LFInst_7_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_7_LFInst_0_U3  ( .A(PermutationOutput[28]), .ZN(
        \SubCellInst_LFInst_7_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_7_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_7_LFInst_1_n5 ), .ZN(Output[29]) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U5  ( .A1(PermutationOutput[30]), 
        .A2(PermutationOutput[28]), .ZN(\SubCellInst_LFInst_7_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_7_LFInst_1_U4  ( .A1(PermutationOutput[31]), .A2(
        \SubCellInst_LFInst_7_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_1_U3  ( .A1(PermutationOutput[30]), 
        .A2(PermutationOutput[28]), .ZN(\SubCellInst_LFInst_7_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_7_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_7_LFInst_2_n10 ), .ZN(Output[30]) );
  OR2_X1 \SubCellInst_LFInst_7_LFInst_2_U7  ( .A1(PermutationOutput[28]), .A2(
        PermutationOutput[31]), .ZN(\SubCellInst_LFInst_7_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U6  ( .A1(PermutationOutput[29]), 
        .A2(\SubCellInst_LFInst_7_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_7_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_7_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U4  ( .A1(PermutationOutput[28]), 
        .A2(PermutationOutput[31]), .ZN(\SubCellInst_LFInst_7_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_7_LFInst_2_U3  ( .A(PermutationOutput[30]), .ZN(
        \SubCellInst_LFInst_7_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_7_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_7_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_7_LFInst_3_n5 ), .ZN(Output[31]) );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_3_U5  ( .A1(PermutationOutput[31]), 
        .A2(PermutationOutput[28]), .ZN(\SubCellInst_LFInst_7_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_3_U4  ( .A1(PermutationOutput[29]), 
        .A2(\SubCellInst_LFInst_7_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_7_LFInst_3_U3  ( .A1(PermutationOutput[31]), 
        .A2(PermutationOutput[30]), .ZN(\SubCellInst_LFInst_7_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_8_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_8_LFInst_0_n10 ), .ZN(Output[32]) );
  AND2_X1 \SubCellInst_LFInst_8_LFInst_0_U7  ( .A1(PermutationOutput[35]), 
        .A2(PermutationOutput[34]), .ZN(\SubCellInst_LFInst_8_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_0_U6  ( .A1(PermutationOutput[33]), 
        .A2(\SubCellInst_LFInst_8_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_8_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_8_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_0_U4  ( .A1(PermutationOutput[35]), 
        .A2(PermutationOutput[34]), .ZN(\SubCellInst_LFInst_8_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_8_LFInst_0_U3  ( .A(PermutationOutput[32]), .ZN(
        \SubCellInst_LFInst_8_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_8_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_8_LFInst_1_n5 ), .ZN(Output[33]) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_1_U5  ( .A1(PermutationOutput[34]), 
        .A2(PermutationOutput[32]), .ZN(\SubCellInst_LFInst_8_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_8_LFInst_1_U4  ( .A1(PermutationOutput[35]), .A2(
        \SubCellInst_LFInst_8_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_1_U3  ( .A1(PermutationOutput[34]), 
        .A2(PermutationOutput[32]), .ZN(\SubCellInst_LFInst_8_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_8_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_8_LFInst_2_n10 ), .ZN(Output[34]) );
  OR2_X1 \SubCellInst_LFInst_8_LFInst_2_U7  ( .A1(PermutationOutput[32]), .A2(
        PermutationOutput[35]), .ZN(\SubCellInst_LFInst_8_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U6  ( .A1(PermutationOutput[33]), 
        .A2(\SubCellInst_LFInst_8_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_8_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_8_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U4  ( .A1(PermutationOutput[32]), 
        .A2(PermutationOutput[35]), .ZN(\SubCellInst_LFInst_8_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_8_LFInst_2_U3  ( .A(PermutationOutput[34]), .ZN(
        \SubCellInst_LFInst_8_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_8_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_8_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_8_LFInst_3_n5 ), .ZN(Output[35]) );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_3_U5  ( .A1(PermutationOutput[35]), 
        .A2(PermutationOutput[32]), .ZN(\SubCellInst_LFInst_8_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_3_U4  ( .A1(PermutationOutput[33]), 
        .A2(\SubCellInst_LFInst_8_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_8_LFInst_3_U3  ( .A1(PermutationOutput[35]), 
        .A2(PermutationOutput[34]), .ZN(\SubCellInst_LFInst_8_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_9_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_9_LFInst_0_n10 ), .ZN(Output[36]) );
  AND2_X1 \SubCellInst_LFInst_9_LFInst_0_U7  ( .A1(PermutationOutput[39]), 
        .A2(PermutationOutput[38]), .ZN(\SubCellInst_LFInst_9_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_0_U6  ( .A1(PermutationOutput[37]), 
        .A2(\SubCellInst_LFInst_9_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_9_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_9_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_0_U4  ( .A1(PermutationOutput[39]), 
        .A2(PermutationOutput[38]), .ZN(\SubCellInst_LFInst_9_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_9_LFInst_0_U3  ( .A(PermutationOutput[36]), .ZN(
        \SubCellInst_LFInst_9_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_9_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_9_LFInst_1_n5 ), .ZN(Output[37]) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_1_U5  ( .A1(PermutationOutput[38]), 
        .A2(PermutationOutput[36]), .ZN(\SubCellInst_LFInst_9_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_9_LFInst_1_U4  ( .A1(PermutationOutput[39]), .A2(
        \SubCellInst_LFInst_9_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_1_U3  ( .A1(PermutationOutput[38]), 
        .A2(PermutationOutput[36]), .ZN(\SubCellInst_LFInst_9_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_9_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_9_LFInst_2_n10 ), .ZN(Output[38]) );
  OR2_X1 \SubCellInst_LFInst_9_LFInst_2_U7  ( .A1(PermutationOutput[36]), .A2(
        PermutationOutput[39]), .ZN(\SubCellInst_LFInst_9_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U6  ( .A1(PermutationOutput[37]), 
        .A2(\SubCellInst_LFInst_9_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_9_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_9_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U4  ( .A1(PermutationOutput[36]), 
        .A2(PermutationOutput[39]), .ZN(\SubCellInst_LFInst_9_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_9_LFInst_2_U3  ( .A(PermutationOutput[38]), .ZN(
        \SubCellInst_LFInst_9_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_9_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_9_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_9_LFInst_3_n5 ), .ZN(Output[39]) );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_3_U5  ( .A1(PermutationOutput[39]), 
        .A2(PermutationOutput[36]), .ZN(\SubCellInst_LFInst_9_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_3_U4  ( .A1(PermutationOutput[37]), 
        .A2(\SubCellInst_LFInst_9_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_9_LFInst_3_U3  ( .A1(PermutationOutput[39]), 
        .A2(PermutationOutput[38]), .ZN(\SubCellInst_LFInst_9_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_10_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_10_LFInst_0_n10 ), .ZN(Output[40]) );
  AND2_X1 \SubCellInst_LFInst_10_LFInst_0_U7  ( .A1(PermutationOutput[43]), 
        .A2(PermutationOutput[42]), .ZN(\SubCellInst_LFInst_10_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_0_U6  ( .A1(PermutationOutput[41]), 
        .A2(\SubCellInst_LFInst_10_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_10_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_10_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_0_U4  ( .A1(PermutationOutput[43]), 
        .A2(PermutationOutput[42]), .ZN(\SubCellInst_LFInst_10_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst_LFInst_10_LFInst_0_U3  ( .A(PermutationOutput[40]), .ZN(
        \SubCellInst_LFInst_10_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_10_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_10_LFInst_1_n5 ), .ZN(Output[41]) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_1_U5  ( .A1(PermutationOutput[42]), 
        .A2(PermutationOutput[40]), .ZN(\SubCellInst_LFInst_10_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst_LFInst_10_LFInst_1_U4  ( .A1(PermutationOutput[43]), 
        .A2(\SubCellInst_LFInst_10_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_1_U3  ( .A1(PermutationOutput[42]), 
        .A2(PermutationOutput[40]), .ZN(\SubCellInst_LFInst_10_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_10_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_10_LFInst_2_n10 ), .ZN(Output[42]) );
  OR2_X1 \SubCellInst_LFInst_10_LFInst_2_U7  ( .A1(PermutationOutput[40]), 
        .A2(PermutationOutput[43]), .ZN(\SubCellInst_LFInst_10_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U6  ( .A1(PermutationOutput[41]), 
        .A2(\SubCellInst_LFInst_10_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_10_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_10_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U4  ( .A1(PermutationOutput[40]), 
        .A2(PermutationOutput[43]), .ZN(\SubCellInst_LFInst_10_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst_LFInst_10_LFInst_2_U3  ( .A(PermutationOutput[42]), .ZN(
        \SubCellInst_LFInst_10_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_10_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_10_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_10_LFInst_3_n5 ), .ZN(Output[43]) );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_3_U5  ( .A1(PermutationOutput[43]), 
        .A2(PermutationOutput[40]), .ZN(\SubCellInst_LFInst_10_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_3_U4  ( .A1(PermutationOutput[41]), 
        .A2(\SubCellInst_LFInst_10_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_10_LFInst_3_U3  ( .A1(PermutationOutput[43]), 
        .A2(PermutationOutput[42]), .ZN(\SubCellInst_LFInst_10_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_11_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_11_LFInst_0_n10 ), .ZN(Output[44]) );
  AND2_X1 \SubCellInst_LFInst_11_LFInst_0_U7  ( .A1(PermutationOutput[47]), 
        .A2(PermutationOutput[46]), .ZN(\SubCellInst_LFInst_11_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_0_U6  ( .A1(PermutationOutput[45]), 
        .A2(\SubCellInst_LFInst_11_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_11_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_11_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_0_U4  ( .A1(PermutationOutput[47]), 
        .A2(PermutationOutput[46]), .ZN(\SubCellInst_LFInst_11_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst_LFInst_11_LFInst_0_U3  ( .A(PermutationOutput[44]), .ZN(
        \SubCellInst_LFInst_11_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_11_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_11_LFInst_1_n5 ), .ZN(Output[45]) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_1_U5  ( .A1(PermutationOutput[46]), 
        .A2(PermutationOutput[44]), .ZN(\SubCellInst_LFInst_11_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst_LFInst_11_LFInst_1_U4  ( .A1(PermutationOutput[47]), 
        .A2(\SubCellInst_LFInst_11_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_1_U3  ( .A1(PermutationOutput[46]), 
        .A2(PermutationOutput[44]), .ZN(\SubCellInst_LFInst_11_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_11_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_11_LFInst_2_n10 ), .ZN(Output[46]) );
  OR2_X1 \SubCellInst_LFInst_11_LFInst_2_U7  ( .A1(PermutationOutput[44]), 
        .A2(PermutationOutput[47]), .ZN(\SubCellInst_LFInst_11_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U6  ( .A1(PermutationOutput[45]), 
        .A2(\SubCellInst_LFInst_11_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_11_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_11_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U4  ( .A1(PermutationOutput[44]), 
        .A2(PermutationOutput[47]), .ZN(\SubCellInst_LFInst_11_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst_LFInst_11_LFInst_2_U3  ( .A(PermutationOutput[46]), .ZN(
        \SubCellInst_LFInst_11_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_11_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_11_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_11_LFInst_3_n5 ), .ZN(Output[47]) );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_3_U5  ( .A1(PermutationOutput[47]), 
        .A2(PermutationOutput[44]), .ZN(\SubCellInst_LFInst_11_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_3_U4  ( .A1(PermutationOutput[45]), 
        .A2(\SubCellInst_LFInst_11_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_11_LFInst_3_U3  ( .A1(PermutationOutput[47]), 
        .A2(PermutationOutput[46]), .ZN(\SubCellInst_LFInst_11_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_12_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_12_LFInst_0_n10 ), .ZN(Output[48]) );
  AND2_X1 \SubCellInst_LFInst_12_LFInst_0_U7  ( .A1(PermutationOutput[51]), 
        .A2(PermutationOutput[50]), .ZN(\SubCellInst_LFInst_12_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_0_U6  ( .A1(PermutationOutput[49]), 
        .A2(\SubCellInst_LFInst_12_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_12_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_12_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_0_U4  ( .A1(PermutationOutput[51]), 
        .A2(PermutationOutput[50]), .ZN(\SubCellInst_LFInst_12_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst_LFInst_12_LFInst_0_U3  ( .A(PermutationOutput[48]), .ZN(
        \SubCellInst_LFInst_12_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_12_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_12_LFInst_1_n5 ), .ZN(Output[49]) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U5  ( .A1(PermutationOutput[50]), 
        .A2(PermutationOutput[48]), .ZN(\SubCellInst_LFInst_12_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst_LFInst_12_LFInst_1_U4  ( .A1(PermutationOutput[51]), 
        .A2(\SubCellInst_LFInst_12_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_1_U3  ( .A1(PermutationOutput[50]), 
        .A2(PermutationOutput[48]), .ZN(\SubCellInst_LFInst_12_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_12_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_12_LFInst_2_n10 ), .ZN(Output[50]) );
  OR2_X1 \SubCellInst_LFInst_12_LFInst_2_U7  ( .A1(PermutationOutput[48]), 
        .A2(PermutationOutput[51]), .ZN(\SubCellInst_LFInst_12_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U6  ( .A1(PermutationOutput[49]), 
        .A2(\SubCellInst_LFInst_12_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_12_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_12_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U4  ( .A1(PermutationOutput[48]), 
        .A2(PermutationOutput[51]), .ZN(\SubCellInst_LFInst_12_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst_LFInst_12_LFInst_2_U3  ( .A(PermutationOutput[50]), .ZN(
        \SubCellInst_LFInst_12_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_12_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_12_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_12_LFInst_3_n5 ), .ZN(Output[51]) );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_3_U5  ( .A1(PermutationOutput[51]), 
        .A2(PermutationOutput[48]), .ZN(\SubCellInst_LFInst_12_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_3_U4  ( .A1(PermutationOutput[49]), 
        .A2(\SubCellInst_LFInst_12_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_12_LFInst_3_U3  ( .A1(PermutationOutput[51]), 
        .A2(PermutationOutput[50]), .ZN(\SubCellInst_LFInst_12_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_13_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_13_LFInst_0_n10 ), .ZN(Output[52]) );
  AND2_X1 \SubCellInst_LFInst_13_LFInst_0_U7  ( .A1(PermutationOutput[55]), 
        .A2(PermutationOutput[54]), .ZN(\SubCellInst_LFInst_13_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_0_U6  ( .A1(PermutationOutput[53]), 
        .A2(\SubCellInst_LFInst_13_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_13_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_13_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_0_U4  ( .A1(PermutationOutput[55]), 
        .A2(PermutationOutput[54]), .ZN(\SubCellInst_LFInst_13_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst_LFInst_13_LFInst_0_U3  ( .A(PermutationOutput[52]), .ZN(
        \SubCellInst_LFInst_13_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_13_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_13_LFInst_1_n5 ), .ZN(Output[53]) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U5  ( .A1(PermutationOutput[54]), 
        .A2(PermutationOutput[52]), .ZN(\SubCellInst_LFInst_13_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst_LFInst_13_LFInst_1_U4  ( .A1(PermutationOutput[55]), 
        .A2(\SubCellInst_LFInst_13_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_1_U3  ( .A1(PermutationOutput[54]), 
        .A2(PermutationOutput[52]), .ZN(\SubCellInst_LFInst_13_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_13_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_13_LFInst_2_n10 ), .ZN(Output[54]) );
  OR2_X1 \SubCellInst_LFInst_13_LFInst_2_U7  ( .A1(PermutationOutput[52]), 
        .A2(PermutationOutput[55]), .ZN(\SubCellInst_LFInst_13_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U6  ( .A1(PermutationOutput[53]), 
        .A2(\SubCellInst_LFInst_13_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_13_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_13_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U4  ( .A1(PermutationOutput[52]), 
        .A2(PermutationOutput[55]), .ZN(\SubCellInst_LFInst_13_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst_LFInst_13_LFInst_2_U3  ( .A(PermutationOutput[54]), .ZN(
        \SubCellInst_LFInst_13_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_13_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_13_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_13_LFInst_3_n5 ), .ZN(Output[55]) );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_3_U5  ( .A1(PermutationOutput[55]), 
        .A2(PermutationOutput[52]), .ZN(\SubCellInst_LFInst_13_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_3_U4  ( .A1(PermutationOutput[53]), 
        .A2(\SubCellInst_LFInst_13_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_13_LFInst_3_U3  ( .A1(PermutationOutput[55]), 
        .A2(PermutationOutput[54]), .ZN(\SubCellInst_LFInst_13_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_14_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_14_LFInst_0_n10 ), .ZN(Output[56]) );
  AND2_X1 \SubCellInst_LFInst_14_LFInst_0_U7  ( .A1(PermutationOutput[59]), 
        .A2(PermutationOutput[58]), .ZN(\SubCellInst_LFInst_14_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_0_U6  ( .A1(PermutationOutput[57]), 
        .A2(\SubCellInst_LFInst_14_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_14_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_14_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_0_U4  ( .A1(PermutationOutput[59]), 
        .A2(PermutationOutput[58]), .ZN(\SubCellInst_LFInst_14_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst_LFInst_14_LFInst_0_U3  ( .A(PermutationOutput[56]), .ZN(
        \SubCellInst_LFInst_14_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_14_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_14_LFInst_1_n5 ), .ZN(Output[57]) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U5  ( .A1(PermutationOutput[58]), 
        .A2(PermutationOutput[56]), .ZN(\SubCellInst_LFInst_14_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst_LFInst_14_LFInst_1_U4  ( .A1(PermutationOutput[59]), 
        .A2(\SubCellInst_LFInst_14_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_1_U3  ( .A1(PermutationOutput[58]), 
        .A2(PermutationOutput[56]), .ZN(\SubCellInst_LFInst_14_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_14_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_14_LFInst_2_n10 ), .ZN(Output[58]) );
  OR2_X1 \SubCellInst_LFInst_14_LFInst_2_U7  ( .A1(PermutationOutput[56]), 
        .A2(PermutationOutput[59]), .ZN(\SubCellInst_LFInst_14_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U6  ( .A1(PermutationOutput[57]), 
        .A2(\SubCellInst_LFInst_14_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_14_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_14_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U4  ( .A1(PermutationOutput[56]), 
        .A2(PermutationOutput[59]), .ZN(\SubCellInst_LFInst_14_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst_LFInst_14_LFInst_2_U3  ( .A(PermutationOutput[58]), .ZN(
        \SubCellInst_LFInst_14_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_14_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_14_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_14_LFInst_3_n5 ), .ZN(Output[59]) );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_3_U5  ( .A1(PermutationOutput[59]), 
        .A2(PermutationOutput[56]), .ZN(\SubCellInst_LFInst_14_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_3_U4  ( .A1(PermutationOutput[57]), 
        .A2(\SubCellInst_LFInst_14_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_14_LFInst_3_U3  ( .A1(PermutationOutput[59]), 
        .A2(PermutationOutput[58]), .ZN(\SubCellInst_LFInst_14_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_15_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_15_LFInst_0_n10 ), .ZN(Output[60]) );
  AND2_X1 \SubCellInst_LFInst_15_LFInst_0_U7  ( .A1(PermutationOutput[63]), 
        .A2(PermutationOutput[62]), .ZN(\SubCellInst_LFInst_15_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_0_U6  ( .A1(PermutationOutput[61]), 
        .A2(\SubCellInst_LFInst_15_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_15_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_15_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_0_U4  ( .A1(PermutationOutput[63]), 
        .A2(PermutationOutput[62]), .ZN(\SubCellInst_LFInst_15_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst_LFInst_15_LFInst_0_U3  ( .A(PermutationOutput[60]), .ZN(
        \SubCellInst_LFInst_15_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_15_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_15_LFInst_1_n5 ), .ZN(Output[61]) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U5  ( .A1(PermutationOutput[62]), 
        .A2(PermutationOutput[60]), .ZN(\SubCellInst_LFInst_15_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst_LFInst_15_LFInst_1_U4  ( .A1(PermutationOutput[63]), 
        .A2(\SubCellInst_LFInst_15_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_1_U3  ( .A1(PermutationOutput[62]), 
        .A2(PermutationOutput[60]), .ZN(\SubCellInst_LFInst_15_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_15_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_15_LFInst_2_n10 ), .ZN(Output[62]) );
  OR2_X1 \SubCellInst_LFInst_15_LFInst_2_U7  ( .A1(PermutationOutput[60]), 
        .A2(PermutationOutput[63]), .ZN(\SubCellInst_LFInst_15_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U6  ( .A1(PermutationOutput[61]), 
        .A2(\SubCellInst_LFInst_15_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_15_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_15_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U4  ( .A1(PermutationOutput[60]), 
        .A2(PermutationOutput[63]), .ZN(\SubCellInst_LFInst_15_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst_LFInst_15_LFInst_2_U3  ( .A(PermutationOutput[62]), .ZN(
        \SubCellInst_LFInst_15_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_15_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_15_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_15_LFInst_3_n5 ), .ZN(Output[63]) );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_3_U5  ( .A1(PermutationOutput[63]), 
        .A2(PermutationOutput[60]), .ZN(\SubCellInst_LFInst_15_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_3_U4  ( .A1(PermutationOutput[61]), 
        .A2(\SubCellInst_LFInst_15_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_15_LFInst_3_U3  ( .A1(PermutationOutput[63]), 
        .A2(PermutationOutput[62]), .ZN(\SubCellInst_LFInst_15_LFInst_3_n4 )
         );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_0_LFInst_0_n2 ), .B(Input[2]), .ZN(
        Red_MCOutput[0]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_0_U3  ( .A(Input[3]), .B(
        Input[1]), .ZN(\Red_PlaintextInst_LFInst_0_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_0_LFInst_1_n2 ), .B(Input[2]), .ZN(
        Red_MCOutput[1]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_1_U3  ( .A(Input[3]), .B(
        Input[0]), .ZN(\Red_PlaintextInst_LFInst_0_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_0_LFInst_2_n2 ), .B(Input[1]), .ZN(
        Red_MCOutput[2]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_2_U3  ( .A(Input[3]), .B(
        Input[0]), .ZN(\Red_PlaintextInst_LFInst_0_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_0_LFInst_3_n2 ), .B(Input[1]), .ZN(
        Red_MCOutput[3]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_3_U3  ( .A(Input[2]), .B(
        Input[0]), .ZN(\Red_PlaintextInst_LFInst_0_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_1_LFInst_0_n2 ), .B(Input[6]), .ZN(
        Red_MCOutput[4]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_0_U3  ( .A(Input[7]), .B(
        Input[5]), .ZN(\Red_PlaintextInst_LFInst_1_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_1_LFInst_1_n2 ), .B(Input[6]), .ZN(
        Red_MCOutput[5]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_1_U3  ( .A(Input[7]), .B(
        Input[4]), .ZN(\Red_PlaintextInst_LFInst_1_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_1_LFInst_2_n2 ), .B(Input[5]), .ZN(
        Red_MCOutput[6]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_2_U3  ( .A(Input[7]), .B(
        Input[4]), .ZN(\Red_PlaintextInst_LFInst_1_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_1_LFInst_3_n2 ), .B(Input[5]), .ZN(
        Red_MCOutput[7]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_3_U3  ( .A(Input[6]), .B(
        Input[4]), .ZN(\Red_PlaintextInst_LFInst_1_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_2_LFInst_0_n2 ), .B(Input[10]), .ZN(
        Red_MCOutput[8]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_0_U3  ( .A(Input[11]), .B(
        Input[9]), .ZN(\Red_PlaintextInst_LFInst_2_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_2_LFInst_1_n2 ), .B(Input[10]), .ZN(
        Red_MCOutput[9]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_1_U3  ( .A(Input[11]), .B(
        Input[8]), .ZN(\Red_PlaintextInst_LFInst_2_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_2_LFInst_2_n2 ), .B(Input[9]), .ZN(
        Red_MCOutput[10]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_2_U3  ( .A(Input[11]), .B(
        Input[8]), .ZN(\Red_PlaintextInst_LFInst_2_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_2_LFInst_3_n2 ), .B(Input[9]), .ZN(
        Red_MCOutput[11]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_3_U3  ( .A(Input[10]), .B(
        Input[8]), .ZN(\Red_PlaintextInst_LFInst_2_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_3_LFInst_0_n2 ), .B(Input[14]), .ZN(
        Red_MCOutput[12]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_0_U3  ( .A(Input[15]), .B(
        Input[13]), .ZN(\Red_PlaintextInst_LFInst_3_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_3_LFInst_1_n2 ), .B(Input[14]), .ZN(
        Red_MCOutput[13]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_1_U3  ( .A(Input[15]), .B(
        Input[12]), .ZN(\Red_PlaintextInst_LFInst_3_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_3_LFInst_2_n2 ), .B(Input[13]), .ZN(
        Red_MCOutput[14]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_2_U3  ( .A(Input[15]), .B(
        Input[12]), .ZN(\Red_PlaintextInst_LFInst_3_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_3_LFInst_3_n2 ), .B(Input[13]), .ZN(
        Red_MCOutput[15]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_3_U3  ( .A(Input[14]), .B(
        Input[12]), .ZN(\Red_PlaintextInst_LFInst_3_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_4_LFInst_0_n2 ), .B(Input[18]), .ZN(
        Red_MCOutput[16]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_0_U3  ( .A(Input[19]), .B(
        Input[17]), .ZN(\Red_PlaintextInst_LFInst_4_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_4_LFInst_1_n2 ), .B(Input[18]), .ZN(
        Red_MCOutput[17]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_1_U3  ( .A(Input[19]), .B(
        Input[16]), .ZN(\Red_PlaintextInst_LFInst_4_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_4_LFInst_2_n2 ), .B(Input[17]), .ZN(
        Red_MCOutput[18]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_2_U3  ( .A(Input[19]), .B(
        Input[16]), .ZN(\Red_PlaintextInst_LFInst_4_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_4_LFInst_3_n2 ), .B(Input[17]), .ZN(
        Red_MCOutput[19]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_3_U3  ( .A(Input[18]), .B(
        Input[16]), .ZN(\Red_PlaintextInst_LFInst_4_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_5_LFInst_0_n2 ), .B(Input[22]), .ZN(
        Red_MCOutput[20]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_0_U3  ( .A(Input[23]), .B(
        Input[21]), .ZN(\Red_PlaintextInst_LFInst_5_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_5_LFInst_1_n2 ), .B(Input[22]), .ZN(
        Red_MCOutput[21]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_1_U3  ( .A(Input[23]), .B(
        Input[20]), .ZN(\Red_PlaintextInst_LFInst_5_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_5_LFInst_2_n2 ), .B(Input[21]), .ZN(
        Red_MCOutput[22]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_2_U3  ( .A(Input[23]), .B(
        Input[20]), .ZN(\Red_PlaintextInst_LFInst_5_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_5_LFInst_3_n2 ), .B(Input[21]), .ZN(
        Red_MCOutput[23]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_3_U3  ( .A(Input[22]), .B(
        Input[20]), .ZN(\Red_PlaintextInst_LFInst_5_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_6_LFInst_0_n2 ), .B(Input[26]), .ZN(
        Red_MCOutput[24]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_0_U3  ( .A(Input[27]), .B(
        Input[25]), .ZN(\Red_PlaintextInst_LFInst_6_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_6_LFInst_1_n2 ), .B(Input[26]), .ZN(
        Red_MCOutput[25]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_1_U3  ( .A(Input[27]), .B(
        Input[24]), .ZN(\Red_PlaintextInst_LFInst_6_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_6_LFInst_2_n2 ), .B(Input[25]), .ZN(
        Red_MCOutput[26]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_2_U3  ( .A(Input[27]), .B(
        Input[24]), .ZN(\Red_PlaintextInst_LFInst_6_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_6_LFInst_3_n2 ), .B(Input[25]), .ZN(
        Red_MCOutput[27]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_3_U3  ( .A(Input[26]), .B(
        Input[24]), .ZN(\Red_PlaintextInst_LFInst_6_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_7_LFInst_0_n2 ), .B(Input[30]), .ZN(
        Red_MCOutput[28]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_0_U3  ( .A(Input[31]), .B(
        Input[29]), .ZN(\Red_PlaintextInst_LFInst_7_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_7_LFInst_1_n2 ), .B(Input[30]), .ZN(
        Red_MCOutput[29]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_1_U3  ( .A(Input[31]), .B(
        Input[28]), .ZN(\Red_PlaintextInst_LFInst_7_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_7_LFInst_2_n2 ), .B(Input[29]), .ZN(
        Red_MCOutput[30]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_2_U3  ( .A(Input[31]), .B(
        Input[28]), .ZN(\Red_PlaintextInst_LFInst_7_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_7_LFInst_3_n2 ), .B(Input[29]), .ZN(
        Red_MCOutput[31]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_3_U3  ( .A(Input[30]), .B(
        Input[28]), .ZN(\Red_PlaintextInst_LFInst_7_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_8_LFInst_0_n2 ), .B(Input[34]), .ZN(
        Red_Input[32]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_0_U3  ( .A(Input[35]), .B(
        Input[33]), .ZN(\Red_PlaintextInst_LFInst_8_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_8_LFInst_1_n2 ), .B(Input[34]), .ZN(
        Red_Input[33]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_1_U3  ( .A(Input[35]), .B(
        Input[32]), .ZN(\Red_PlaintextInst_LFInst_8_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_8_LFInst_2_n2 ), .B(Input[33]), .ZN(
        Red_Input[34]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_2_U3  ( .A(Input[35]), .B(
        Input[32]), .ZN(\Red_PlaintextInst_LFInst_8_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_8_LFInst_3_n2 ), .B(Input[33]), .ZN(
        Red_Input[35]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_3_U3  ( .A(Input[34]), .B(
        Input[32]), .ZN(\Red_PlaintextInst_LFInst_8_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_9_LFInst_0_n2 ), .B(Input[38]), .ZN(
        Red_Input[36]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_0_U3  ( .A(Input[39]), .B(
        Input[37]), .ZN(\Red_PlaintextInst_LFInst_9_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_9_LFInst_1_n2 ), .B(Input[38]), .ZN(
        Red_Input[37]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_1_U3  ( .A(Input[39]), .B(
        Input[36]), .ZN(\Red_PlaintextInst_LFInst_9_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_9_LFInst_2_n2 ), .B(Input[37]), .ZN(
        Red_Input[38]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_2_U3  ( .A(Input[39]), .B(
        Input[36]), .ZN(\Red_PlaintextInst_LFInst_9_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_9_LFInst_3_n2 ), .B(Input[37]), .ZN(
        Red_Input[39]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_3_U3  ( .A(Input[38]), .B(
        Input[36]), .ZN(\Red_PlaintextInst_LFInst_9_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_10_LFInst_0_n2 ), .B(Input[42]), .ZN(
        Red_Input[40]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_0_U3  ( .A(Input[43]), .B(
        Input[41]), .ZN(\Red_PlaintextInst_LFInst_10_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_10_LFInst_1_n2 ), .B(Input[42]), .ZN(
        Red_Input[41]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_1_U3  ( .A(Input[43]), .B(
        Input[40]), .ZN(\Red_PlaintextInst_LFInst_10_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_10_LFInst_2_n2 ), .B(Input[41]), .ZN(
        Red_Input[42]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_2_U3  ( .A(Input[43]), .B(
        Input[40]), .ZN(\Red_PlaintextInst_LFInst_10_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_10_LFInst_3_n2 ), .B(Input[41]), .ZN(
        Red_Input[43]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_3_U3  ( .A(Input[42]), .B(
        Input[40]), .ZN(\Red_PlaintextInst_LFInst_10_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_11_LFInst_0_n2 ), .B(Input[46]), .ZN(
        Red_Input[44]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_0_U3  ( .A(Input[47]), .B(
        Input[45]), .ZN(\Red_PlaintextInst_LFInst_11_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_11_LFInst_1_n2 ), .B(Input[46]), .ZN(
        Red_Input[45]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_1_U3  ( .A(Input[47]), .B(
        Input[44]), .ZN(\Red_PlaintextInst_LFInst_11_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_11_LFInst_2_n2 ), .B(Input[45]), .ZN(
        Red_Input[46]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_2_U3  ( .A(Input[47]), .B(
        Input[44]), .ZN(\Red_PlaintextInst_LFInst_11_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_11_LFInst_3_n2 ), .B(Input[45]), .ZN(
        Red_Input[47]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_3_U3  ( .A(Input[46]), .B(
        Input[44]), .ZN(\Red_PlaintextInst_LFInst_11_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_12_LFInst_0_n2 ), .B(Input[50]), .ZN(
        Red_Input[48]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_0_U3  ( .A(Input[51]), .B(
        Input[49]), .ZN(\Red_PlaintextInst_LFInst_12_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_12_LFInst_1_n2 ), .B(Input[50]), .ZN(
        Red_Input[49]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_1_U3  ( .A(Input[51]), .B(
        Input[48]), .ZN(\Red_PlaintextInst_LFInst_12_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_12_LFInst_2_n2 ), .B(Input[49]), .ZN(
        Red_Input[50]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_2_U3  ( .A(Input[51]), .B(
        Input[48]), .ZN(\Red_PlaintextInst_LFInst_12_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_12_LFInst_3_n2 ), .B(Input[49]), .ZN(
        Red_Input[51]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_3_U3  ( .A(Input[50]), .B(
        Input[48]), .ZN(\Red_PlaintextInst_LFInst_12_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_13_LFInst_0_n2 ), .B(Input[54]), .ZN(
        Red_Input[52]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_0_U3  ( .A(Input[55]), .B(
        Input[53]), .ZN(\Red_PlaintextInst_LFInst_13_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_13_LFInst_1_n2 ), .B(Input[54]), .ZN(
        Red_Input[53]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_1_U3  ( .A(Input[55]), .B(
        Input[52]), .ZN(\Red_PlaintextInst_LFInst_13_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_13_LFInst_2_n2 ), .B(Input[53]), .ZN(
        Red_Input[54]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_2_U3  ( .A(Input[55]), .B(
        Input[52]), .ZN(\Red_PlaintextInst_LFInst_13_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_13_LFInst_3_n2 ), .B(Input[53]), .ZN(
        Red_Input[55]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_3_U3  ( .A(Input[54]), .B(
        Input[52]), .ZN(\Red_PlaintextInst_LFInst_13_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_14_LFInst_0_n2 ), .B(Input[58]), .ZN(
        Red_Input[56]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_0_U3  ( .A(Input[59]), .B(
        Input[57]), .ZN(\Red_PlaintextInst_LFInst_14_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_14_LFInst_1_n2 ), .B(Input[58]), .ZN(
        Red_Input[57]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_1_U3  ( .A(Input[59]), .B(
        Input[56]), .ZN(\Red_PlaintextInst_LFInst_14_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_14_LFInst_2_n2 ), .B(Input[57]), .ZN(
        Red_Input[58]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_2_U3  ( .A(Input[59]), .B(
        Input[56]), .ZN(\Red_PlaintextInst_LFInst_14_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_14_LFInst_3_n2 ), .B(Input[57]), .ZN(
        Red_Input[59]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_3_U3  ( .A(Input[58]), .B(
        Input[56]), .ZN(\Red_PlaintextInst_LFInst_14_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_15_LFInst_0_n2 ), .B(Input[62]), .ZN(
        Red_Input[60]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_0_U3  ( .A(Input[63]), .B(
        Input[61]), .ZN(\Red_PlaintextInst_LFInst_15_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_15_LFInst_1_n2 ), .B(Input[62]), .ZN(
        Red_Input[61]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_1_U3  ( .A(Input[63]), .B(
        Input[60]), .ZN(\Red_PlaintextInst_LFInst_15_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_15_LFInst_2_n2 ), .B(Input[61]), .ZN(
        Red_Input[62]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_2_U3  ( .A(Input[63]), .B(
        Input[60]), .ZN(\Red_PlaintextInst_LFInst_15_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_15_LFInst_3_n2 ), .B(Input[61]), .ZN(
        Red_Input[63]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_3_U3  ( .A(Input[62]), .B(
        Input[60]), .ZN(\Red_PlaintextInst_LFInst_15_LFInst_3_n2 ) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_0_U2  ( .A(\Red_MCInst_XOR_r0_Inst_0_n3 ), 
        .B(Red_MCOutput[0]), .ZN(Red_MCOutput[48]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_0_U1  ( .A(Red_Input[48]), .B(
        Red_MCOutput[16]), .ZN(\Red_MCInst_XOR_r0_Inst_0_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_0_U1  ( .A(Red_Input[32]), .B(
        Red_MCOutput[0]), .Z(Red_MCOutput[32]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_1_U2  ( .A(\Red_MCInst_XOR_r0_Inst_1_n3 ), 
        .B(Red_MCOutput[1]), .ZN(Red_MCOutput[49]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_1_U1  ( .A(Red_Input[49]), .B(
        Red_MCOutput[17]), .ZN(\Red_MCInst_XOR_r0_Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_1_U1  ( .A(Red_Input[33]), .B(
        Red_MCOutput[1]), .Z(Red_MCOutput[33]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_2_U2  ( .A(\Red_MCInst_XOR_r0_Inst_2_n3 ), 
        .B(Red_MCOutput[2]), .ZN(Red_MCOutput[50]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_2_U1  ( .A(Red_Input[50]), .B(
        Red_MCOutput[18]), .ZN(\Red_MCInst_XOR_r0_Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_2_U1  ( .A(Red_Input[34]), .B(
        Red_MCOutput[2]), .Z(Red_MCOutput[34]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_3_U2  ( .A(\Red_MCInst_XOR_r0_Inst_3_n3 ), 
        .B(Red_MCOutput[3]), .ZN(Red_MCOutput[51]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_3_U1  ( .A(Red_Input[51]), .B(
        Red_MCOutput[19]), .ZN(\Red_MCInst_XOR_r0_Inst_3_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_3_U1  ( .A(Red_Input[35]), .B(
        Red_MCOutput[3]), .Z(Red_MCOutput[35]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_4_U2  ( .A(\Red_MCInst_XOR_r0_Inst_4_n3 ), 
        .B(Red_MCOutput[4]), .ZN(Red_MCOutput[52]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_4_U1  ( .A(Red_Input[52]), .B(
        Red_MCOutput[20]), .ZN(\Red_MCInst_XOR_r0_Inst_4_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_4_U1  ( .A(Red_Input[36]), .B(
        Red_MCOutput[4]), .Z(Red_MCOutput[36]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_5_U2  ( .A(\Red_MCInst_XOR_r0_Inst_5_n3 ), 
        .B(Red_MCOutput[5]), .ZN(Red_MCOutput[53]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_5_U1  ( .A(Red_Input[53]), .B(
        Red_MCOutput[21]), .ZN(\Red_MCInst_XOR_r0_Inst_5_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_5_U1  ( .A(Red_Input[37]), .B(
        Red_MCOutput[5]), .Z(Red_MCOutput[37]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_6_U2  ( .A(\Red_MCInst_XOR_r0_Inst_6_n3 ), 
        .B(Red_MCOutput[6]), .ZN(Red_MCOutput[54]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_6_U1  ( .A(Red_Input[54]), .B(
        Red_MCOutput[22]), .ZN(\Red_MCInst_XOR_r0_Inst_6_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_6_U1  ( .A(Red_Input[38]), .B(
        Red_MCOutput[6]), .Z(Red_MCOutput[38]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_7_U2  ( .A(\Red_MCInst_XOR_r0_Inst_7_n3 ), 
        .B(Red_MCOutput[7]), .ZN(Red_MCOutput[55]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_7_U1  ( .A(Red_Input[55]), .B(
        Red_MCOutput[23]), .ZN(\Red_MCInst_XOR_r0_Inst_7_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_7_U1  ( .A(Red_Input[39]), .B(
        Red_MCOutput[7]), .Z(Red_MCOutput[39]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_8_U2  ( .A(\Red_MCInst_XOR_r0_Inst_8_n3 ), 
        .B(Red_MCOutput[8]), .ZN(Red_MCOutput[56]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_8_U1  ( .A(Red_Input[56]), .B(
        Red_MCOutput[24]), .ZN(\Red_MCInst_XOR_r0_Inst_8_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_8_U1  ( .A(Red_Input[40]), .B(
        Red_MCOutput[8]), .Z(Red_MCOutput[40]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_9_U2  ( .A(\Red_MCInst_XOR_r0_Inst_9_n3 ), 
        .B(Red_MCOutput[9]), .ZN(Red_MCOutput[57]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_9_U1  ( .A(Red_Input[57]), .B(
        Red_MCOutput[25]), .ZN(\Red_MCInst_XOR_r0_Inst_9_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_9_U1  ( .A(Red_Input[41]), .B(
        Red_MCOutput[9]), .Z(Red_MCOutput[41]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_10_U2  ( .A(\Red_MCInst_XOR_r0_Inst_10_n3 ), 
        .B(Red_MCOutput[10]), .ZN(Red_MCOutput[58]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_10_U1  ( .A(Red_Input[58]), .B(
        Red_MCOutput[26]), .ZN(\Red_MCInst_XOR_r0_Inst_10_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_10_U1  ( .A(Red_Input[42]), .B(
        Red_MCOutput[10]), .Z(Red_MCOutput[42]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_11_U2  ( .A(\Red_MCInst_XOR_r0_Inst_11_n3 ), 
        .B(Red_MCOutput[11]), .ZN(Red_MCOutput[59]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_11_U1  ( .A(Red_Input[59]), .B(
        Red_MCOutput[27]), .ZN(\Red_MCInst_XOR_r0_Inst_11_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_11_U1  ( .A(Red_Input[43]), .B(
        Red_MCOutput[11]), .Z(Red_MCOutput[43]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_12_U2  ( .A(\Red_MCInst_XOR_r0_Inst_12_n3 ), 
        .B(Red_MCOutput[12]), .ZN(Red_MCOutput[60]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_12_U1  ( .A(Red_Input[60]), .B(
        Red_MCOutput[28]), .ZN(\Red_MCInst_XOR_r0_Inst_12_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_12_U1  ( .A(Red_Input[44]), .B(
        Red_MCOutput[12]), .Z(Red_MCOutput[44]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_13_U2  ( .A(\Red_MCInst_XOR_r0_Inst_13_n3 ), 
        .B(Red_MCOutput[13]), .ZN(Red_MCOutput[61]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_13_U1  ( .A(Red_Input[61]), .B(
        Red_MCOutput[29]), .ZN(\Red_MCInst_XOR_r0_Inst_13_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_13_U1  ( .A(Red_Input[45]), .B(
        Red_MCOutput[13]), .Z(Red_MCOutput[45]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_14_U2  ( .A(\Red_MCInst_XOR_r0_Inst_14_n3 ), 
        .B(Red_MCOutput[14]), .ZN(Red_MCOutput[62]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_14_U1  ( .A(Red_Input[62]), .B(
        Red_MCOutput[30]), .ZN(\Red_MCInst_XOR_r0_Inst_14_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_14_U1  ( .A(Red_Input[46]), .B(
        Red_MCOutput[14]), .Z(Red_MCOutput[46]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_15_U2  ( .A(\Red_MCInst_XOR_r0_Inst_15_n3 ), 
        .B(Red_MCOutput[15]), .ZN(Red_MCOutput[63]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_15_U1  ( .A(Red_Input[63]), .B(
        Red_MCOutput[31]), .ZN(\Red_MCInst_XOR_r0_Inst_15_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_15_U1  ( .A(Red_Input[47]), .B(
        Red_MCOutput[15]), .Z(Red_MCOutput[47]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_0_0_U1  ( .A(Red_MCOutput[48]), .B(
        Red_K0[48]), .Z(Red_AddRoundKeyOutput[48]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_0_1_U1  ( .A(Red_MCOutput[49]), .B(
        Red_K0[49]), .Z(Red_AddRoundKeyOutput[49]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_0_2_U1  ( .A(Red_MCOutput[50]), .B(
        Red_K0[50]), .Z(Red_AddRoundKeyOutput[50]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_0_3_U1  ( .A(Red_MCOutput[51]), .B(
        Red_K0[51]), .Z(Red_AddRoundKeyOutput[51]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_1_0_U1  ( .A(Red_MCOutput[52]), .B(
        Red_K0[52]), .Z(Red_AddRoundKeyOutput[52]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_1_1_U1  ( .A(Red_MCOutput[53]), .B(
        Red_K0[53]), .Z(Red_AddRoundKeyOutput[53]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_1_2_U1  ( .A(Red_MCOutput[54]), .B(
        Red_K0[54]), .Z(Red_AddRoundKeyOutput[54]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_1_3_U1  ( .A(Red_MCOutput[55]), .B(
        Red_K0[55]), .Z(Red_AddRoundKeyOutput[55]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_2_0_U1  ( .A(Red_MCOutput[56]), .B(
        Red_K0[56]), .Z(Red_AddRoundKeyOutput[56]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_2_1_U1  ( .A(Red_MCOutput[57]), .B(
        Red_K0[57]), .Z(Red_AddRoundKeyOutput[57]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_2_2_U1  ( .A(Red_MCOutput[58]), .B(
        Red_K0[58]), .Z(Red_AddRoundKeyOutput[58]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_2_3_U1  ( .A(Red_MCOutput[59]), .B(
        Red_K0[59]), .Z(Red_AddRoundKeyOutput[59]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_3_0_U1  ( .A(Red_MCOutput[60]), .B(
        Red_K0[60]), .Z(Red_AddRoundKeyOutput[60]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_3_1_U1  ( .A(Red_MCOutput[61]), .B(
        Red_K0[61]), .Z(Red_AddRoundKeyOutput[61]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_3_2_U1  ( .A(Red_MCOutput[62]), .B(
        Red_K0[62]), .Z(Red_AddRoundKeyOutput[62]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_3_3_U1  ( .A(Red_MCOutput[63]), .B(
        Red_K0[63]), .Z(Red_AddRoundKeyOutput[63]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_0_0_U1  ( .A(Red_K0[40]), .B(
        Red_MCOutput[40]), .Z(Red_AddRoundKeyOutput[40]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_0_1_U1  ( .A(Red_K0[41]), .B(
        Red_MCOutput[41]), .Z(Red_AddRoundKeyOutput[41]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_0_2_U1  ( .A(Red_K0[42]), .B(
        Red_MCOutput[42]), .Z(Red_AddRoundKeyOutput[42]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_0_3_U1  ( .A(Red_K0[43]), .B(
        Red_MCOutput[43]), .Z(Red_AddRoundKeyOutput[43]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_1_0_U1  ( .A(Red_K0[44]), .B(
        Red_MCOutput[44]), .Z(Red_AddRoundKeyOutput[44]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_1_1_U1  ( .A(Red_K0[45]), .B(
        Red_MCOutput[45]), .Z(Red_AddRoundKeyOutput[45]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_1_2_U1  ( .A(Red_K0[46]), .B(
        Red_MCOutput[46]), .Z(Red_AddRoundKeyOutput[46]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_1_3_U1  ( .A(Red_K0[47]), .B(
        Red_MCOutput[47]), .Z(Red_AddRoundKeyOutput[47]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_0_0_U1  ( .A(Red_MCOutput[0]), .B(Red_K0[0]), 
        .Z(Red_AddRoundKeyOutput[0]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_0_1_U1  ( .A(Red_MCOutput[1]), .B(Red_K0[1]), 
        .Z(Red_AddRoundKeyOutput[1]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_0_2_U1  ( .A(Red_MCOutput[2]), .B(Red_K0[2]), 
        .Z(Red_AddRoundKeyOutput[2]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_0_3_U1  ( .A(Red_MCOutput[3]), .B(Red_K0[3]), 
        .Z(Red_AddRoundKeyOutput[3]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_1_0_U1  ( .A(Red_MCOutput[4]), .B(Red_K0[4]), 
        .Z(Red_AddRoundKeyOutput[4]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_1_1_U1  ( .A(Red_MCOutput[5]), .B(Red_K0[5]), 
        .Z(Red_AddRoundKeyOutput[5]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_1_2_U1  ( .A(Red_MCOutput[6]), .B(Red_K0[6]), 
        .Z(Red_AddRoundKeyOutput[6]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_1_3_U1  ( .A(Red_MCOutput[7]), .B(Red_K0[7]), 
        .Z(Red_AddRoundKeyOutput[7]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_2_0_U1  ( .A(Red_MCOutput[8]), .B(Red_K0[8]), 
        .Z(Red_AddRoundKeyOutput[8]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_2_1_U1  ( .A(Red_MCOutput[9]), .B(Red_K0[9]), 
        .Z(Red_AddRoundKeyOutput[9]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_2_2_U1  ( .A(Red_MCOutput[10]), .B(
        Red_K0[10]), .Z(Red_AddRoundKeyOutput[10]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_2_3_U1  ( .A(Red_MCOutput[11]), .B(
        Red_K0[11]), .Z(Red_AddRoundKeyOutput[11]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_3_0_U1  ( .A(Red_MCOutput[12]), .B(
        Red_K0[12]), .Z(Red_AddRoundKeyOutput[12]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_3_1_U1  ( .A(Red_MCOutput[13]), .B(
        Red_K0[13]), .Z(Red_AddRoundKeyOutput[13]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_3_2_U1  ( .A(Red_MCOutput[14]), .B(
        Red_K0[14]), .Z(Red_AddRoundKeyOutput[14]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_3_3_U1  ( .A(Red_MCOutput[15]), .B(
        Red_K0[15]), .Z(Red_AddRoundKeyOutput[15]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_4_0_U1  ( .A(Red_MCOutput[16]), .B(
        Red_K0[16]), .Z(Red_AddRoundKeyOutput[16]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_4_1_U1  ( .A(Red_MCOutput[17]), .B(
        Red_K0[17]), .Z(Red_AddRoundKeyOutput[17]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_4_2_U1  ( .A(Red_MCOutput[18]), .B(
        Red_K0[18]), .Z(Red_AddRoundKeyOutput[18]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_4_3_U1  ( .A(Red_MCOutput[19]), .B(
        Red_K0[19]), .Z(Red_AddRoundKeyOutput[19]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_5_0_U1  ( .A(Red_MCOutput[20]), .B(
        Red_K0[20]), .Z(Red_AddRoundKeyOutput[20]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_5_1_U1  ( .A(Red_MCOutput[21]), .B(
        Red_K0[21]), .Z(Red_AddRoundKeyOutput[21]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_5_2_U1  ( .A(Red_MCOutput[22]), .B(
        Red_K0[22]), .Z(Red_AddRoundKeyOutput[22]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_5_3_U1  ( .A(Red_MCOutput[23]), .B(
        Red_K0[23]), .Z(Red_AddRoundKeyOutput[23]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_6_0_U1  ( .A(Red_MCOutput[24]), .B(
        Red_K0[24]), .Z(Red_AddRoundKeyOutput[24]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_6_1_U1  ( .A(Red_MCOutput[25]), .B(
        Red_K0[25]), .Z(Red_AddRoundKeyOutput[25]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_6_2_U1  ( .A(Red_MCOutput[26]), .B(
        Red_K0[26]), .Z(Red_AddRoundKeyOutput[26]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_6_3_U1  ( .A(Red_MCOutput[27]), .B(
        Red_K0[27]), .Z(Red_AddRoundKeyOutput[27]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_7_0_U1  ( .A(Red_MCOutput[28]), .B(
        Red_K0[28]), .Z(Red_AddRoundKeyOutput[28]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_7_1_U1  ( .A(Red_MCOutput[29]), .B(
        Red_K0[29]), .Z(Red_AddRoundKeyOutput[29]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_7_2_U1  ( .A(Red_MCOutput[30]), .B(
        Red_K0[30]), .Z(Red_AddRoundKeyOutput[30]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_7_3_U1  ( .A(Red_MCOutput[31]), .B(
        Red_K0[31]), .Z(Red_AddRoundKeyOutput[31]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_8_0_U1  ( .A(Red_MCOutput[32]), .B(
        Red_K0[32]), .Z(Red_AddRoundKeyOutput[32]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_8_1_U1  ( .A(Red_MCOutput[33]), .B(
        Red_K0[33]), .Z(Red_AddRoundKeyOutput[33]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_8_2_U1  ( .A(Red_MCOutput[34]), .B(
        Red_K0[34]), .Z(Red_AddRoundKeyOutput[34]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_8_3_U1  ( .A(Red_MCOutput[35]), .B(
        Red_K0[35]), .Z(Red_AddRoundKeyOutput[35]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_9_0_U1  ( .A(Red_MCOutput[36]), .B(
        Red_K0[36]), .Z(Red_AddRoundKeyOutput[36]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_9_1_U1  ( .A(Red_MCOutput[37]), .B(
        Red_K0[37]), .Z(Red_AddRoundKeyOutput[37]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_9_2_U1  ( .A(Red_MCOutput[38]), .B(
        Red_K0[38]), .Z(Red_AddRoundKeyOutput[38]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_9_3_U1  ( .A(Red_MCOutput[39]), .B(
        Red_K0[39]), .Z(Red_AddRoundKeyOutput[39]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[0]  ( .D(Red_AddRoundKeyOutput[0]), 
        .CK(clk), .Q(Red_StateRegOutput[0]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[1]  ( .D(Red_AddRoundKeyOutput[1]), 
        .CK(clk), .Q(Red_StateRegOutput[1]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[2]  ( .D(Red_AddRoundKeyOutput[2]), 
        .CK(clk), .Q(Red_StateRegOutput[2]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[3]  ( .D(Red_AddRoundKeyOutput[3]), 
        .CK(clk), .Q(Red_StateRegOutput[3]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[4]  ( .D(Red_AddRoundKeyOutput[4]), 
        .CK(clk), .Q(Red_StateRegOutput[4]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[5]  ( .D(Red_AddRoundKeyOutput[5]), 
        .CK(clk), .Q(Red_StateRegOutput[5]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[6]  ( .D(Red_AddRoundKeyOutput[6]), 
        .CK(clk), .Q(Red_StateRegOutput[6]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[7]  ( .D(Red_AddRoundKeyOutput[7]), 
        .CK(clk), .Q(Red_StateRegOutput[7]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[8]  ( .D(Red_AddRoundKeyOutput[8]), 
        .CK(clk), .Q(Red_StateRegOutput[8]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[9]  ( .D(Red_AddRoundKeyOutput[9]), 
        .CK(clk), .Q(Red_StateRegOutput[9]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[10]  ( .D(Red_AddRoundKeyOutput[10]), .CK(clk), .Q(Red_StateRegOutput[10]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[11]  ( .D(Red_AddRoundKeyOutput[11]), .CK(clk), .Q(Red_StateRegOutput[11]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[12]  ( .D(Red_AddRoundKeyOutput[12]), .CK(clk), .Q(Red_StateRegOutput[12]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[13]  ( .D(Red_AddRoundKeyOutput[13]), .CK(clk), .Q(Red_StateRegOutput[13]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[14]  ( .D(Red_AddRoundKeyOutput[14]), .CK(clk), .Q(Red_StateRegOutput[14]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[15]  ( .D(Red_AddRoundKeyOutput[15]), .CK(clk), .Q(Red_StateRegOutput[15]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[16]  ( .D(Red_AddRoundKeyOutput[16]), .CK(clk), .Q(Red_StateRegOutput[16]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[17]  ( .D(Red_AddRoundKeyOutput[17]), .CK(clk), .Q(Red_StateRegOutput[17]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[18]  ( .D(Red_AddRoundKeyOutput[18]), .CK(clk), .Q(Red_StateRegOutput[18]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[19]  ( .D(Red_AddRoundKeyOutput[19]), .CK(clk), .Q(Red_StateRegOutput[19]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[20]  ( .D(Red_AddRoundKeyOutput[20]), .CK(clk), .Q(Red_StateRegOutput[20]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[21]  ( .D(Red_AddRoundKeyOutput[21]), .CK(clk), .Q(Red_StateRegOutput[21]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[22]  ( .D(Red_AddRoundKeyOutput[22]), .CK(clk), .Q(Red_StateRegOutput[22]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[23]  ( .D(Red_AddRoundKeyOutput[23]), .CK(clk), .Q(Red_StateRegOutput[23]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[24]  ( .D(Red_AddRoundKeyOutput[24]), .CK(clk), .Q(Red_StateRegOutput[24]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[25]  ( .D(Red_AddRoundKeyOutput[25]), .CK(clk), .Q(Red_StateRegOutput[25]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[26]  ( .D(Red_AddRoundKeyOutput[26]), .CK(clk), .Q(Red_StateRegOutput[26]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[27]  ( .D(Red_AddRoundKeyOutput[27]), .CK(clk), .Q(Red_StateRegOutput[27]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[28]  ( .D(Red_AddRoundKeyOutput[28]), .CK(clk), .Q(Red_StateRegOutput[28]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[29]  ( .D(Red_AddRoundKeyOutput[29]), .CK(clk), .Q(Red_StateRegOutput[29]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[30]  ( .D(Red_AddRoundKeyOutput[30]), .CK(clk), .Q(Red_StateRegOutput[30]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[31]  ( .D(Red_AddRoundKeyOutput[31]), .CK(clk), .Q(Red_StateRegOutput[31]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[32]  ( .D(Red_AddRoundKeyOutput[32]), .CK(clk), .Q(Red_StateRegOutput[32]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[33]  ( .D(Red_AddRoundKeyOutput[33]), .CK(clk), .Q(Red_StateRegOutput[33]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[34]  ( .D(Red_AddRoundKeyOutput[34]), .CK(clk), .Q(Red_StateRegOutput[34]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[35]  ( .D(Red_AddRoundKeyOutput[35]), .CK(clk), .Q(Red_StateRegOutput[35]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[36]  ( .D(Red_AddRoundKeyOutput[36]), .CK(clk), .Q(Red_StateRegOutput[36]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[37]  ( .D(Red_AddRoundKeyOutput[37]), .CK(clk), .Q(Red_StateRegOutput[37]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[38]  ( .D(Red_AddRoundKeyOutput[38]), .CK(clk), .Q(Red_StateRegOutput[38]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[39]  ( .D(Red_AddRoundKeyOutput[39]), .CK(clk), .Q(Red_StateRegOutput[39]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[40]  ( .D(Red_AddRoundKeyOutput[40]), .CK(clk), .Q(Red_StateRegOutput[40]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[41]  ( .D(Red_AddRoundKeyOutput[41]), .CK(clk), .Q(Red_StateRegOutput[41]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[42]  ( .D(Red_AddRoundKeyOutput[42]), .CK(clk), .Q(Red_StateRegOutput[42]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[43]  ( .D(Red_AddRoundKeyOutput[43]), .CK(clk), .Q(Red_StateRegOutput[43]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[44]  ( .D(Red_AddRoundKeyOutput[44]), .CK(clk), .Q(Red_StateRegOutput[44]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[45]  ( .D(Red_AddRoundKeyOutput[45]), .CK(clk), .Q(Red_StateRegOutput[45]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[46]  ( .D(Red_AddRoundKeyOutput[46]), .CK(clk), .Q(Red_StateRegOutput[46]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[47]  ( .D(Red_AddRoundKeyOutput[47]), .CK(clk), .Q(Red_StateRegOutput[47]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[48]  ( .D(Red_AddRoundKeyOutput[48]), .CK(clk), .Q(Red_StateRegOutput[48]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[49]  ( .D(Red_AddRoundKeyOutput[49]), .CK(clk), .Q(Red_StateRegOutput[49]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[50]  ( .D(Red_AddRoundKeyOutput[50]), .CK(clk), .Q(Red_StateRegOutput[50]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[51]  ( .D(Red_AddRoundKeyOutput[51]), .CK(clk), .Q(Red_StateRegOutput[51]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[52]  ( .D(Red_AddRoundKeyOutput[52]), .CK(clk), .Q(Red_StateRegOutput[52]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[53]  ( .D(Red_AddRoundKeyOutput[53]), .CK(clk), .Q(Red_StateRegOutput[53]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[54]  ( .D(Red_AddRoundKeyOutput[54]), .CK(clk), .Q(Red_StateRegOutput[54]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[55]  ( .D(Red_AddRoundKeyOutput[55]), .CK(clk), .Q(Red_StateRegOutput[55]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[56]  ( .D(Red_AddRoundKeyOutput[56]), .CK(clk), .Q(Red_StateRegOutput[56]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[57]  ( .D(Red_AddRoundKeyOutput[57]), .CK(clk), .Q(Red_StateRegOutput[57]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[58]  ( .D(Red_AddRoundKeyOutput[58]), .CK(clk), .Q(Red_StateRegOutput[58]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[59]  ( .D(Red_AddRoundKeyOutput[59]), .CK(clk), .Q(Red_StateRegOutput[59]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[60]  ( .D(Red_AddRoundKeyOutput[60]), .CK(clk), .Q(Red_StateRegOutput[60]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[61]  ( .D(Red_AddRoundKeyOutput[61]), .CK(clk), .Q(Red_StateRegOutput[61]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[62]  ( .D(Red_AddRoundKeyOutput[62]), .CK(clk), .Q(Red_StateRegOutput[62]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[63]  ( .D(Red_AddRoundKeyOutput[63]), .CK(clk), .Q(Red_StateRegOutput[63]) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_0_LFInst_0_n13 ), .ZN(Red_Feedback[0]) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U9  ( .A1(PermutationOutput[0]), 
        .A2(\Red_SubCellInst_LFInst_0_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_0_n11 ), .A2(PermutationOutput[2]), 
        .ZN(\Red_SubCellInst_LFInst_0_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_0_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_0_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U6  ( .A1(PermutationOutput[3]), 
        .A2(\Red_SubCellInst_LFInst_0_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U5  ( .A(PermutationOutput[1]), 
        .ZN(\Red_SubCellInst_LFInst_0_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U4  ( .A1(PermutationOutput[2]), 
        .A2(\Red_SubCellInst_LFInst_0_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U3  ( .A(PermutationOutput[0]), 
        .ZN(\Red_SubCellInst_LFInst_0_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_0_LFInst_1_n14 ), .ZN(Red_Feedback[1]) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_1_n13 ), .A2(PermutationOutput[1]), 
        .ZN(\Red_SubCellInst_LFInst_0_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_1_n12 ), .A2(PermutationOutput[0]), 
        .ZN(\Red_SubCellInst_LFInst_0_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_1_U5  ( .A1(PermutationOutput[3]), 
        .A2(PermutationOutput[2]), .ZN(\Red_SubCellInst_LFInst_0_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_0_LFInst_1_U4  ( .A1(PermutationOutput[2]), 
        .A2(\Red_SubCellInst_LFInst_0_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_1_U3  ( .A(PermutationOutput[0]), 
        .B(PermutationOutput[3]), .ZN(\Red_SubCellInst_LFInst_0_LFInst_1_n11 )
         );
  NOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_0_LFInst_2_n18 ), .ZN(Red_Feedback[2]) );
  AND2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_2_n17 ), .A2(PermutationOutput[0]), 
        .ZN(\Red_SubCellInst_LFInst_0_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U8  ( .A1(PermutationOutput[2]), 
        .A2(PermutationOutput[1]), .ZN(\Red_SubCellInst_LFInst_0_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_0_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_0_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U6  ( .A1(PermutationOutput[3]), 
        .A2(\Red_SubCellInst_LFInst_0_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U5  ( .A(PermutationOutput[1]), 
        .ZN(\Red_SubCellInst_LFInst_0_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U4  ( .A1(PermutationOutput[2]), 
        .A2(\Red_SubCellInst_LFInst_0_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U3  ( .A(PermutationOutput[0]), 
        .ZN(\Red_SubCellInst_LFInst_0_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_3_U6  ( .A(PermutationOutput[1]), 
        .B(\Red_SubCellInst_LFInst_0_LFInst_3_n8 ), .ZN(Red_Feedback[3]) );
  NOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_0_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_3_U4  ( .A1(PermutationOutput[2]), 
        .A2(PermutationOutput[3]), .ZN(\Red_SubCellInst_LFInst_0_LFInst_3_n6 )
         );
  AND2_X1 \Red_SubCellInst_LFInst_0_LFInst_3_U3  ( .A1(PermutationOutput[3]), 
        .A2(PermutationOutput[0]), .ZN(\Red_SubCellInst_LFInst_0_LFInst_3_n7 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_1_LFInst_0_n13 ), .ZN(Red_Feedback[4]) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U9  ( .A1(PermutationOutput[4]), 
        .A2(\Red_SubCellInst_LFInst_1_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_0_n11 ), .A2(PermutationOutput[6]), 
        .ZN(\Red_SubCellInst_LFInst_1_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_1_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_1_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U6  ( .A1(PermutationOutput[7]), 
        .A2(\Red_SubCellInst_LFInst_1_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U5  ( .A(PermutationOutput[5]), 
        .ZN(\Red_SubCellInst_LFInst_1_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U4  ( .A1(PermutationOutput[6]), 
        .A2(\Red_SubCellInst_LFInst_1_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U3  ( .A(PermutationOutput[4]), 
        .ZN(\Red_SubCellInst_LFInst_1_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_1_LFInst_1_n14 ), .ZN(Red_Feedback[5]) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_1_n13 ), .A2(PermutationOutput[5]), 
        .ZN(\Red_SubCellInst_LFInst_1_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_1_n12 ), .A2(PermutationOutput[4]), 
        .ZN(\Red_SubCellInst_LFInst_1_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_1_U5  ( .A1(PermutationOutput[7]), 
        .A2(PermutationOutput[6]), .ZN(\Red_SubCellInst_LFInst_1_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_1_LFInst_1_U4  ( .A1(PermutationOutput[6]), 
        .A2(\Red_SubCellInst_LFInst_1_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_1_U3  ( .A(PermutationOutput[4]), 
        .B(PermutationOutput[7]), .ZN(\Red_SubCellInst_LFInst_1_LFInst_1_n11 )
         );
  NOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_1_LFInst_2_n18 ), .ZN(Red_Feedback[6]) );
  AND2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_2_n17 ), .A2(PermutationOutput[4]), 
        .ZN(\Red_SubCellInst_LFInst_1_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U8  ( .A1(PermutationOutput[6]), 
        .A2(PermutationOutput[5]), .ZN(\Red_SubCellInst_LFInst_1_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_1_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_1_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U6  ( .A1(PermutationOutput[7]), 
        .A2(\Red_SubCellInst_LFInst_1_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U5  ( .A(PermutationOutput[5]), 
        .ZN(\Red_SubCellInst_LFInst_1_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U4  ( .A1(PermutationOutput[6]), 
        .A2(\Red_SubCellInst_LFInst_1_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U3  ( .A(PermutationOutput[4]), 
        .ZN(\Red_SubCellInst_LFInst_1_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_3_U6  ( .A(PermutationOutput[5]), 
        .B(\Red_SubCellInst_LFInst_1_LFInst_3_n8 ), .ZN(Red_Feedback[7]) );
  NOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_1_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_3_U4  ( .A1(PermutationOutput[6]), 
        .A2(PermutationOutput[7]), .ZN(\Red_SubCellInst_LFInst_1_LFInst_3_n6 )
         );
  AND2_X1 \Red_SubCellInst_LFInst_1_LFInst_3_U3  ( .A1(PermutationOutput[7]), 
        .A2(PermutationOutput[4]), .ZN(\Red_SubCellInst_LFInst_1_LFInst_3_n7 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_2_LFInst_0_n13 ), .ZN(Red_Feedback[8]) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U9  ( .A1(PermutationOutput[8]), 
        .A2(\Red_SubCellInst_LFInst_2_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_0_n11 ), .A2(PermutationOutput[10]), 
        .ZN(\Red_SubCellInst_LFInst_2_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_2_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_2_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U6  ( .A1(PermutationOutput[11]), 
        .A2(\Red_SubCellInst_LFInst_2_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U5  ( .A(PermutationOutput[9]), 
        .ZN(\Red_SubCellInst_LFInst_2_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U4  ( .A1(PermutationOutput[10]), 
        .A2(\Red_SubCellInst_LFInst_2_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U3  ( .A(PermutationOutput[8]), 
        .ZN(\Red_SubCellInst_LFInst_2_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_2_LFInst_1_n14 ), .ZN(Red_Feedback[9]) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_1_n13 ), .A2(PermutationOutput[9]), 
        .ZN(\Red_SubCellInst_LFInst_2_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_1_n12 ), .A2(PermutationOutput[8]), 
        .ZN(\Red_SubCellInst_LFInst_2_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_1_U5  ( .A1(PermutationOutput[11]), 
        .A2(PermutationOutput[10]), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_2_LFInst_1_U4  ( .A1(PermutationOutput[10]), 
        .A2(\Red_SubCellInst_LFInst_2_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_1_U3  ( .A(PermutationOutput[8]), 
        .B(PermutationOutput[11]), .ZN(\Red_SubCellInst_LFInst_2_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_2_LFInst_2_n18 ), .ZN(Red_Feedback[10]) );
  AND2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_2_n17 ), .A2(PermutationOutput[8]), 
        .ZN(\Red_SubCellInst_LFInst_2_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U8  ( .A1(PermutationOutput[10]), 
        .A2(PermutationOutput[9]), .ZN(\Red_SubCellInst_LFInst_2_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_2_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_2_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U6  ( .A1(PermutationOutput[11]), 
        .A2(\Red_SubCellInst_LFInst_2_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U5  ( .A(PermutationOutput[9]), 
        .ZN(\Red_SubCellInst_LFInst_2_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U4  ( .A1(PermutationOutput[10]), 
        .A2(\Red_SubCellInst_LFInst_2_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U3  ( .A(PermutationOutput[8]), 
        .ZN(\Red_SubCellInst_LFInst_2_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_3_U6  ( .A(PermutationOutput[9]), 
        .B(\Red_SubCellInst_LFInst_2_LFInst_3_n8 ), .ZN(Red_Feedback[11]) );
  NOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_2_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_3_U4  ( .A1(PermutationOutput[10]), 
        .A2(PermutationOutput[11]), .ZN(\Red_SubCellInst_LFInst_2_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_2_LFInst_3_U3  ( .A1(PermutationOutput[11]), 
        .A2(PermutationOutput[8]), .ZN(\Red_SubCellInst_LFInst_2_LFInst_3_n7 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_3_LFInst_0_n13 ), .ZN(Red_Feedback[12]) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U9  ( .A1(PermutationOutput[12]), 
        .A2(\Red_SubCellInst_LFInst_3_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_0_n11 ), .A2(PermutationOutput[14]), 
        .ZN(\Red_SubCellInst_LFInst_3_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_3_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_3_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U6  ( .A1(PermutationOutput[15]), 
        .A2(\Red_SubCellInst_LFInst_3_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U5  ( .A(PermutationOutput[13]), 
        .ZN(\Red_SubCellInst_LFInst_3_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U4  ( .A1(PermutationOutput[14]), 
        .A2(\Red_SubCellInst_LFInst_3_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U3  ( .A(PermutationOutput[12]), 
        .ZN(\Red_SubCellInst_LFInst_3_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_3_LFInst_1_n14 ), .ZN(Red_Feedback[13]) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_1_n13 ), .A2(PermutationOutput[13]), 
        .ZN(\Red_SubCellInst_LFInst_3_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_1_n12 ), .A2(PermutationOutput[12]), 
        .ZN(\Red_SubCellInst_LFInst_3_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_1_U5  ( .A1(PermutationOutput[15]), 
        .A2(PermutationOutput[14]), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_3_LFInst_1_U4  ( .A1(PermutationOutput[14]), 
        .A2(\Red_SubCellInst_LFInst_3_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_1_U3  ( .A(PermutationOutput[12]), 
        .B(PermutationOutput[15]), .ZN(\Red_SubCellInst_LFInst_3_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_3_LFInst_2_n18 ), .ZN(Red_Feedback[14]) );
  AND2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_2_n17 ), .A2(PermutationOutput[12]), 
        .ZN(\Red_SubCellInst_LFInst_3_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U8  ( .A1(PermutationOutput[14]), 
        .A2(PermutationOutput[13]), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_3_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_3_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U6  ( .A1(PermutationOutput[15]), 
        .A2(\Red_SubCellInst_LFInst_3_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U5  ( .A(PermutationOutput[13]), 
        .ZN(\Red_SubCellInst_LFInst_3_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U4  ( .A1(PermutationOutput[14]), 
        .A2(\Red_SubCellInst_LFInst_3_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U3  ( .A(PermutationOutput[12]), 
        .ZN(\Red_SubCellInst_LFInst_3_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_3_U6  ( .A(PermutationOutput[13]), 
        .B(\Red_SubCellInst_LFInst_3_LFInst_3_n8 ), .ZN(Red_Feedback[15]) );
  NOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_3_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_3_U4  ( .A1(PermutationOutput[14]), 
        .A2(PermutationOutput[15]), .ZN(\Red_SubCellInst_LFInst_3_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_3_LFInst_3_U3  ( .A1(PermutationOutput[15]), 
        .A2(PermutationOutput[12]), .ZN(\Red_SubCellInst_LFInst_3_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_4_LFInst_0_n13 ), .ZN(Red_Feedback[16]) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U9  ( .A1(PermutationOutput[16]), 
        .A2(\Red_SubCellInst_LFInst_4_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_0_n11 ), .A2(PermutationOutput[18]), 
        .ZN(\Red_SubCellInst_LFInst_4_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_4_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_4_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U6  ( .A1(PermutationOutput[19]), 
        .A2(\Red_SubCellInst_LFInst_4_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U5  ( .A(PermutationOutput[17]), 
        .ZN(\Red_SubCellInst_LFInst_4_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U4  ( .A1(PermutationOutput[18]), 
        .A2(\Red_SubCellInst_LFInst_4_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U3  ( .A(PermutationOutput[16]), 
        .ZN(\Red_SubCellInst_LFInst_4_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_4_LFInst_1_n14 ), .ZN(Red_Feedback[17]) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_1_n13 ), .A2(PermutationOutput[17]), 
        .ZN(\Red_SubCellInst_LFInst_4_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_1_n12 ), .A2(PermutationOutput[16]), 
        .ZN(\Red_SubCellInst_LFInst_4_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_1_U5  ( .A1(PermutationOutput[19]), 
        .A2(PermutationOutput[18]), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_4_LFInst_1_U4  ( .A1(PermutationOutput[18]), 
        .A2(\Red_SubCellInst_LFInst_4_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_1_U3  ( .A(PermutationOutput[16]), 
        .B(PermutationOutput[19]), .ZN(\Red_SubCellInst_LFInst_4_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_4_LFInst_2_n18 ), .ZN(Red_Feedback[18]) );
  AND2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_2_n17 ), .A2(PermutationOutput[16]), 
        .ZN(\Red_SubCellInst_LFInst_4_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U8  ( .A1(PermutationOutput[18]), 
        .A2(PermutationOutput[17]), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_4_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_4_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U6  ( .A1(PermutationOutput[19]), 
        .A2(\Red_SubCellInst_LFInst_4_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U5  ( .A(PermutationOutput[17]), 
        .ZN(\Red_SubCellInst_LFInst_4_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U4  ( .A1(PermutationOutput[18]), 
        .A2(\Red_SubCellInst_LFInst_4_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U3  ( .A(PermutationOutput[16]), 
        .ZN(\Red_SubCellInst_LFInst_4_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_3_U6  ( .A(PermutationOutput[17]), 
        .B(\Red_SubCellInst_LFInst_4_LFInst_3_n8 ), .ZN(Red_Feedback[19]) );
  NOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_4_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_3_U4  ( .A1(PermutationOutput[18]), 
        .A2(PermutationOutput[19]), .ZN(\Red_SubCellInst_LFInst_4_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_4_LFInst_3_U3  ( .A1(PermutationOutput[19]), 
        .A2(PermutationOutput[16]), .ZN(\Red_SubCellInst_LFInst_4_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_5_LFInst_0_n13 ), .ZN(Red_Feedback[20]) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U9  ( .A1(PermutationOutput[20]), 
        .A2(\Red_SubCellInst_LFInst_5_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_0_n11 ), .A2(PermutationOutput[22]), 
        .ZN(\Red_SubCellInst_LFInst_5_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_5_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_5_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U6  ( .A1(PermutationOutput[23]), 
        .A2(\Red_SubCellInst_LFInst_5_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U5  ( .A(PermutationOutput[21]), 
        .ZN(\Red_SubCellInst_LFInst_5_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U4  ( .A1(PermutationOutput[22]), 
        .A2(\Red_SubCellInst_LFInst_5_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U3  ( .A(PermutationOutput[20]), 
        .ZN(\Red_SubCellInst_LFInst_5_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_5_LFInst_1_n14 ), .ZN(Red_Feedback[21]) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_1_n13 ), .A2(PermutationOutput[21]), 
        .ZN(\Red_SubCellInst_LFInst_5_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_1_n12 ), .A2(PermutationOutput[20]), 
        .ZN(\Red_SubCellInst_LFInst_5_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_1_U5  ( .A1(PermutationOutput[23]), 
        .A2(PermutationOutput[22]), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_5_LFInst_1_U4  ( .A1(PermutationOutput[22]), 
        .A2(\Red_SubCellInst_LFInst_5_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_1_U3  ( .A(PermutationOutput[20]), 
        .B(PermutationOutput[23]), .ZN(\Red_SubCellInst_LFInst_5_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_5_LFInst_2_n18 ), .ZN(Red_Feedback[22]) );
  AND2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_2_n17 ), .A2(PermutationOutput[20]), 
        .ZN(\Red_SubCellInst_LFInst_5_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U8  ( .A1(PermutationOutput[22]), 
        .A2(PermutationOutput[21]), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_5_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_5_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U6  ( .A1(PermutationOutput[23]), 
        .A2(\Red_SubCellInst_LFInst_5_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U5  ( .A(PermutationOutput[21]), 
        .ZN(\Red_SubCellInst_LFInst_5_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U4  ( .A1(PermutationOutput[22]), 
        .A2(\Red_SubCellInst_LFInst_5_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U3  ( .A(PermutationOutput[20]), 
        .ZN(\Red_SubCellInst_LFInst_5_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_3_U6  ( .A(PermutationOutput[21]), 
        .B(\Red_SubCellInst_LFInst_5_LFInst_3_n8 ), .ZN(Red_Feedback[23]) );
  NOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_5_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_3_U4  ( .A1(PermutationOutput[22]), 
        .A2(PermutationOutput[23]), .ZN(\Red_SubCellInst_LFInst_5_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_5_LFInst_3_U3  ( .A1(PermutationOutput[23]), 
        .A2(PermutationOutput[20]), .ZN(\Red_SubCellInst_LFInst_5_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_6_LFInst_0_n13 ), .ZN(Red_Feedback[24]) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U9  ( .A1(PermutationOutput[24]), 
        .A2(\Red_SubCellInst_LFInst_6_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_0_n11 ), .A2(PermutationOutput[26]), 
        .ZN(\Red_SubCellInst_LFInst_6_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_6_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_6_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U6  ( .A1(PermutationOutput[27]), 
        .A2(\Red_SubCellInst_LFInst_6_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U5  ( .A(PermutationOutput[25]), 
        .ZN(\Red_SubCellInst_LFInst_6_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U4  ( .A1(PermutationOutput[26]), 
        .A2(\Red_SubCellInst_LFInst_6_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U3  ( .A(PermutationOutput[24]), 
        .ZN(\Red_SubCellInst_LFInst_6_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_6_LFInst_1_n14 ), .ZN(Red_Feedback[25]) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_1_n13 ), .A2(PermutationOutput[25]), 
        .ZN(\Red_SubCellInst_LFInst_6_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_1_n12 ), .A2(PermutationOutput[24]), 
        .ZN(\Red_SubCellInst_LFInst_6_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_1_U5  ( .A1(PermutationOutput[27]), 
        .A2(PermutationOutput[26]), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_6_LFInst_1_U4  ( .A1(PermutationOutput[26]), 
        .A2(\Red_SubCellInst_LFInst_6_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_1_U3  ( .A(PermutationOutput[24]), 
        .B(PermutationOutput[27]), .ZN(\Red_SubCellInst_LFInst_6_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_6_LFInst_2_n18 ), .ZN(Red_Feedback[26]) );
  AND2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_2_n17 ), .A2(PermutationOutput[24]), 
        .ZN(\Red_SubCellInst_LFInst_6_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U8  ( .A1(PermutationOutput[26]), 
        .A2(PermutationOutput[25]), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_6_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_6_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U6  ( .A1(PermutationOutput[27]), 
        .A2(\Red_SubCellInst_LFInst_6_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U5  ( .A(PermutationOutput[25]), 
        .ZN(\Red_SubCellInst_LFInst_6_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U4  ( .A1(PermutationOutput[26]), 
        .A2(\Red_SubCellInst_LFInst_6_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U3  ( .A(PermutationOutput[24]), 
        .ZN(\Red_SubCellInst_LFInst_6_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_3_U6  ( .A(PermutationOutput[25]), 
        .B(\Red_SubCellInst_LFInst_6_LFInst_3_n8 ), .ZN(Red_Feedback[27]) );
  NOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_6_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_3_U4  ( .A1(PermutationOutput[26]), 
        .A2(PermutationOutput[27]), .ZN(\Red_SubCellInst_LFInst_6_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_6_LFInst_3_U3  ( .A1(PermutationOutput[27]), 
        .A2(PermutationOutput[24]), .ZN(\Red_SubCellInst_LFInst_6_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_7_LFInst_0_n13 ), .ZN(Red_Feedback[28]) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U9  ( .A1(PermutationOutput[28]), 
        .A2(\Red_SubCellInst_LFInst_7_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_0_n11 ), .A2(PermutationOutput[30]), 
        .ZN(\Red_SubCellInst_LFInst_7_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_7_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_7_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U6  ( .A1(PermutationOutput[31]), 
        .A2(\Red_SubCellInst_LFInst_7_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U5  ( .A(PermutationOutput[29]), 
        .ZN(\Red_SubCellInst_LFInst_7_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U4  ( .A1(PermutationOutput[30]), 
        .A2(\Red_SubCellInst_LFInst_7_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U3  ( .A(PermutationOutput[28]), 
        .ZN(\Red_SubCellInst_LFInst_7_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_7_LFInst_1_n14 ), .ZN(Red_Feedback[29]) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_1_n13 ), .A2(PermutationOutput[29]), 
        .ZN(\Red_SubCellInst_LFInst_7_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_1_n12 ), .A2(PermutationOutput[28]), 
        .ZN(\Red_SubCellInst_LFInst_7_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_1_U5  ( .A1(PermutationOutput[31]), 
        .A2(PermutationOutput[30]), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_7_LFInst_1_U4  ( .A1(PermutationOutput[30]), 
        .A2(\Red_SubCellInst_LFInst_7_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_1_U3  ( .A(PermutationOutput[28]), 
        .B(PermutationOutput[31]), .ZN(\Red_SubCellInst_LFInst_7_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_7_LFInst_2_n18 ), .ZN(Red_Feedback[30]) );
  AND2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_2_n17 ), .A2(PermutationOutput[28]), 
        .ZN(\Red_SubCellInst_LFInst_7_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U8  ( .A1(PermutationOutput[30]), 
        .A2(PermutationOutput[29]), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_7_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_7_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U6  ( .A1(PermutationOutput[31]), 
        .A2(\Red_SubCellInst_LFInst_7_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U5  ( .A(PermutationOutput[29]), 
        .ZN(\Red_SubCellInst_LFInst_7_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U4  ( .A1(PermutationOutput[30]), 
        .A2(\Red_SubCellInst_LFInst_7_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U3  ( .A(PermutationOutput[28]), 
        .ZN(\Red_SubCellInst_LFInst_7_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_3_U6  ( .A(PermutationOutput[29]), 
        .B(\Red_SubCellInst_LFInst_7_LFInst_3_n8 ), .ZN(Red_Feedback[31]) );
  NOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_7_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_3_U4  ( .A1(PermutationOutput[30]), 
        .A2(PermutationOutput[31]), .ZN(\Red_SubCellInst_LFInst_7_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_7_LFInst_3_U3  ( .A1(PermutationOutput[31]), 
        .A2(PermutationOutput[28]), .ZN(\Red_SubCellInst_LFInst_7_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_8_LFInst_0_n13 ), .ZN(Red_Feedback[32]) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U9  ( .A1(PermutationOutput[32]), 
        .A2(\Red_SubCellInst_LFInst_8_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_0_n11 ), .A2(PermutationOutput[34]), 
        .ZN(\Red_SubCellInst_LFInst_8_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_8_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_8_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U6  ( .A1(PermutationOutput[35]), 
        .A2(\Red_SubCellInst_LFInst_8_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U5  ( .A(PermutationOutput[33]), 
        .ZN(\Red_SubCellInst_LFInst_8_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U4  ( .A1(PermutationOutput[34]), 
        .A2(\Red_SubCellInst_LFInst_8_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U3  ( .A(PermutationOutput[32]), 
        .ZN(\Red_SubCellInst_LFInst_8_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_8_LFInst_1_n14 ), .ZN(Red_Feedback[33]) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_1_n13 ), .A2(PermutationOutput[33]), 
        .ZN(\Red_SubCellInst_LFInst_8_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_1_n12 ), .A2(PermutationOutput[32]), 
        .ZN(\Red_SubCellInst_LFInst_8_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_1_U5  ( .A1(PermutationOutput[35]), 
        .A2(PermutationOutput[34]), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_8_LFInst_1_U4  ( .A1(PermutationOutput[34]), 
        .A2(\Red_SubCellInst_LFInst_8_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_1_U3  ( .A(PermutationOutput[32]), 
        .B(PermutationOutput[35]), .ZN(\Red_SubCellInst_LFInst_8_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_8_LFInst_2_n18 ), .ZN(Red_Feedback[34]) );
  AND2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_2_n17 ), .A2(PermutationOutput[32]), 
        .ZN(\Red_SubCellInst_LFInst_8_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U8  ( .A1(PermutationOutput[34]), 
        .A2(PermutationOutput[33]), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_8_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_8_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U6  ( .A1(PermutationOutput[35]), 
        .A2(\Red_SubCellInst_LFInst_8_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U5  ( .A(PermutationOutput[33]), 
        .ZN(\Red_SubCellInst_LFInst_8_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U4  ( .A1(PermutationOutput[34]), 
        .A2(\Red_SubCellInst_LFInst_8_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U3  ( .A(PermutationOutput[32]), 
        .ZN(\Red_SubCellInst_LFInst_8_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_3_U6  ( .A(PermutationOutput[33]), 
        .B(\Red_SubCellInst_LFInst_8_LFInst_3_n8 ), .ZN(Red_Feedback[35]) );
  NOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_8_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_3_U4  ( .A1(PermutationOutput[34]), 
        .A2(PermutationOutput[35]), .ZN(\Red_SubCellInst_LFInst_8_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_8_LFInst_3_U3  ( .A1(PermutationOutput[35]), 
        .A2(PermutationOutput[32]), .ZN(\Red_SubCellInst_LFInst_8_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_9_LFInst_0_n13 ), .ZN(Red_Feedback[36]) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U9  ( .A1(PermutationOutput[36]), 
        .A2(\Red_SubCellInst_LFInst_9_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_0_n11 ), .A2(PermutationOutput[38]), 
        .ZN(\Red_SubCellInst_LFInst_9_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_9_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_9_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U6  ( .A1(PermutationOutput[39]), 
        .A2(\Red_SubCellInst_LFInst_9_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U5  ( .A(PermutationOutput[37]), 
        .ZN(\Red_SubCellInst_LFInst_9_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U4  ( .A1(PermutationOutput[38]), 
        .A2(\Red_SubCellInst_LFInst_9_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U3  ( .A(PermutationOutput[36]), 
        .ZN(\Red_SubCellInst_LFInst_9_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_9_LFInst_1_n14 ), .ZN(Red_Feedback[37]) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_1_n13 ), .A2(PermutationOutput[37]), 
        .ZN(\Red_SubCellInst_LFInst_9_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_1_n12 ), .A2(PermutationOutput[36]), 
        .ZN(\Red_SubCellInst_LFInst_9_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_1_U5  ( .A1(PermutationOutput[39]), 
        .A2(PermutationOutput[38]), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_9_LFInst_1_U4  ( .A1(PermutationOutput[38]), 
        .A2(\Red_SubCellInst_LFInst_9_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_1_U3  ( .A(PermutationOutput[36]), 
        .B(PermutationOutput[39]), .ZN(\Red_SubCellInst_LFInst_9_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_9_LFInst_2_n18 ), .ZN(Red_Feedback[38]) );
  AND2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_2_n17 ), .A2(PermutationOutput[36]), 
        .ZN(\Red_SubCellInst_LFInst_9_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U8  ( .A1(PermutationOutput[38]), 
        .A2(PermutationOutput[37]), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_9_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_9_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U6  ( .A1(PermutationOutput[39]), 
        .A2(\Red_SubCellInst_LFInst_9_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U5  ( .A(PermutationOutput[37]), 
        .ZN(\Red_SubCellInst_LFInst_9_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U4  ( .A1(PermutationOutput[38]), 
        .A2(\Red_SubCellInst_LFInst_9_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U3  ( .A(PermutationOutput[36]), 
        .ZN(\Red_SubCellInst_LFInst_9_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_3_U6  ( .A(PermutationOutput[37]), 
        .B(\Red_SubCellInst_LFInst_9_LFInst_3_n8 ), .ZN(Red_Feedback[39]) );
  NOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_9_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_3_U4  ( .A1(PermutationOutput[38]), 
        .A2(PermutationOutput[39]), .ZN(\Red_SubCellInst_LFInst_9_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_9_LFInst_3_U3  ( .A1(PermutationOutput[39]), 
        .A2(PermutationOutput[36]), .ZN(\Red_SubCellInst_LFInst_9_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_10_LFInst_0_n13 ), .ZN(Red_Feedback[40]) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U9  ( .A1(PermutationOutput[40]), .A2(\Red_SubCellInst_LFInst_10_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_0_n11 ), .A2(PermutationOutput[42]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_10_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_10_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U6  ( .A1(PermutationOutput[43]), .A2(\Red_SubCellInst_LFInst_10_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U5  ( .A(PermutationOutput[41]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U4  ( .A1(PermutationOutput[42]), .A2(\Red_SubCellInst_LFInst_10_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U3  ( .A(PermutationOutput[40]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_10_LFInst_1_n14 ), .ZN(Red_Feedback[41]) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_1_n13 ), .A2(PermutationOutput[41]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_1_n12 ), .A2(PermutationOutput[40]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_1_U5  ( .A1(PermutationOutput[43]), .A2(PermutationOutput[42]), .ZN(\Red_SubCellInst_LFInst_10_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_10_LFInst_1_U4  ( .A1(PermutationOutput[42]), 
        .A2(\Red_SubCellInst_LFInst_10_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_1_U3  ( .A(PermutationOutput[40]), 
        .B(PermutationOutput[43]), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_10_LFInst_2_n18 ), .ZN(Red_Feedback[42]) );
  AND2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_2_n17 ), .A2(PermutationOutput[40]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U8  ( .A1(PermutationOutput[42]), 
        .A2(PermutationOutput[41]), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_10_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_10_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U6  ( .A1(PermutationOutput[43]), 
        .A2(\Red_SubCellInst_LFInst_10_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U5  ( .A(PermutationOutput[41]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U4  ( .A1(PermutationOutput[42]), .A2(\Red_SubCellInst_LFInst_10_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U3  ( .A(PermutationOutput[40]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_3_U6  ( .A(PermutationOutput[41]), 
        .B(\Red_SubCellInst_LFInst_10_LFInst_3_n8 ), .ZN(Red_Feedback[43]) );
  NOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_10_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_3_U4  ( .A1(PermutationOutput[42]), 
        .A2(PermutationOutput[43]), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_10_LFInst_3_U3  ( .A1(PermutationOutput[43]), 
        .A2(PermutationOutput[40]), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_11_LFInst_0_n13 ), .ZN(Red_Feedback[44]) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U9  ( .A1(PermutationOutput[44]), .A2(\Red_SubCellInst_LFInst_11_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_0_n11 ), .A2(PermutationOutput[46]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_11_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_11_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U6  ( .A1(PermutationOutput[47]), .A2(\Red_SubCellInst_LFInst_11_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U5  ( .A(PermutationOutput[45]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U4  ( .A1(PermutationOutput[46]), .A2(\Red_SubCellInst_LFInst_11_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U3  ( .A(PermutationOutput[44]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_11_LFInst_1_n14 ), .ZN(Red_Feedback[45]) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_1_n13 ), .A2(PermutationOutput[45]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_1_n12 ), .A2(PermutationOutput[44]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_1_U5  ( .A1(PermutationOutput[47]), .A2(PermutationOutput[46]), .ZN(\Red_SubCellInst_LFInst_11_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_11_LFInst_1_U4  ( .A1(PermutationOutput[46]), 
        .A2(\Red_SubCellInst_LFInst_11_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_1_U3  ( .A(PermutationOutput[44]), 
        .B(PermutationOutput[47]), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_11_LFInst_2_n18 ), .ZN(Red_Feedback[46]) );
  AND2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_2_n17 ), .A2(PermutationOutput[44]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U8  ( .A1(PermutationOutput[46]), 
        .A2(PermutationOutput[45]), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_11_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_11_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U6  ( .A1(PermutationOutput[47]), 
        .A2(\Red_SubCellInst_LFInst_11_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U5  ( .A(PermutationOutput[45]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U4  ( .A1(PermutationOutput[46]), .A2(\Red_SubCellInst_LFInst_11_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U3  ( .A(PermutationOutput[44]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_3_U6  ( .A(PermutationOutput[45]), 
        .B(\Red_SubCellInst_LFInst_11_LFInst_3_n8 ), .ZN(Red_Feedback[47]) );
  NOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_11_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_3_U4  ( .A1(PermutationOutput[46]), 
        .A2(PermutationOutput[47]), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_11_LFInst_3_U3  ( .A1(PermutationOutput[47]), 
        .A2(PermutationOutput[44]), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_12_LFInst_0_n13 ), .ZN(Red_Feedback[48]) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U9  ( .A1(PermutationOutput[48]), .A2(\Red_SubCellInst_LFInst_12_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_0_n11 ), .A2(PermutationOutput[50]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_12_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_12_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U6  ( .A1(PermutationOutput[51]), .A2(\Red_SubCellInst_LFInst_12_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U5  ( .A(PermutationOutput[49]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U4  ( .A1(PermutationOutput[50]), .A2(\Red_SubCellInst_LFInst_12_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U3  ( .A(PermutationOutput[48]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_12_LFInst_1_n14 ), .ZN(Red_Feedback[49]) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_1_n13 ), .A2(PermutationOutput[49]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_1_n12 ), .A2(PermutationOutput[48]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_1_U5  ( .A1(PermutationOutput[51]), .A2(PermutationOutput[50]), .ZN(\Red_SubCellInst_LFInst_12_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_12_LFInst_1_U4  ( .A1(PermutationOutput[50]), 
        .A2(\Red_SubCellInst_LFInst_12_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_1_U3  ( .A(PermutationOutput[48]), 
        .B(PermutationOutput[51]), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_12_LFInst_2_n18 ), .ZN(Red_Feedback[50]) );
  AND2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_2_n17 ), .A2(PermutationOutput[48]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U8  ( .A1(PermutationOutput[50]), 
        .A2(PermutationOutput[49]), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_12_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_12_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U6  ( .A1(PermutationOutput[51]), 
        .A2(\Red_SubCellInst_LFInst_12_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U5  ( .A(PermutationOutput[49]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U4  ( .A1(PermutationOutput[50]), .A2(\Red_SubCellInst_LFInst_12_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U3  ( .A(PermutationOutput[48]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_3_U6  ( .A(PermutationOutput[49]), 
        .B(\Red_SubCellInst_LFInst_12_LFInst_3_n8 ), .ZN(Red_Feedback[51]) );
  NOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_12_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_3_U4  ( .A1(PermutationOutput[50]), 
        .A2(PermutationOutput[51]), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_12_LFInst_3_U3  ( .A1(PermutationOutput[51]), 
        .A2(PermutationOutput[48]), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_13_LFInst_0_n13 ), .ZN(Red_Feedback[52]) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U9  ( .A1(PermutationOutput[52]), .A2(\Red_SubCellInst_LFInst_13_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_0_n11 ), .A2(PermutationOutput[54]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_13_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_13_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U6  ( .A1(PermutationOutput[55]), .A2(\Red_SubCellInst_LFInst_13_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U5  ( .A(PermutationOutput[53]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U4  ( .A1(PermutationOutput[54]), .A2(\Red_SubCellInst_LFInst_13_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U3  ( .A(PermutationOutput[52]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_13_LFInst_1_n14 ), .ZN(Red_Feedback[53]) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_1_n13 ), .A2(PermutationOutput[53]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_1_n12 ), .A2(PermutationOutput[52]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_1_U5  ( .A1(PermutationOutput[55]), .A2(PermutationOutput[54]), .ZN(\Red_SubCellInst_LFInst_13_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_13_LFInst_1_U4  ( .A1(PermutationOutput[54]), 
        .A2(\Red_SubCellInst_LFInst_13_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_1_U3  ( .A(PermutationOutput[52]), 
        .B(PermutationOutput[55]), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_13_LFInst_2_n18 ), .ZN(Red_Feedback[54]) );
  AND2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_2_n17 ), .A2(PermutationOutput[52]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U8  ( .A1(PermutationOutput[54]), 
        .A2(PermutationOutput[53]), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_13_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_13_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U6  ( .A1(PermutationOutput[55]), 
        .A2(\Red_SubCellInst_LFInst_13_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U5  ( .A(PermutationOutput[53]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U4  ( .A1(PermutationOutput[54]), .A2(\Red_SubCellInst_LFInst_13_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U3  ( .A(PermutationOutput[52]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_3_U6  ( .A(PermutationOutput[53]), 
        .B(\Red_SubCellInst_LFInst_13_LFInst_3_n8 ), .ZN(Red_Feedback[55]) );
  NOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_13_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_3_U4  ( .A1(PermutationOutput[54]), 
        .A2(PermutationOutput[55]), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_13_LFInst_3_U3  ( .A1(PermutationOutput[55]), 
        .A2(PermutationOutput[52]), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_14_LFInst_0_n13 ), .ZN(Red_Feedback[56]) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U9  ( .A1(PermutationOutput[56]), .A2(\Red_SubCellInst_LFInst_14_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_0_n11 ), .A2(PermutationOutput[58]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_14_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_14_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U6  ( .A1(PermutationOutput[59]), .A2(\Red_SubCellInst_LFInst_14_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U5  ( .A(PermutationOutput[57]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U4  ( .A1(PermutationOutput[58]), .A2(\Red_SubCellInst_LFInst_14_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U3  ( .A(PermutationOutput[56]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_14_LFInst_1_n14 ), .ZN(Red_Feedback[57]) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_1_n13 ), .A2(PermutationOutput[57]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_1_n12 ), .A2(PermutationOutput[56]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_1_U5  ( .A1(PermutationOutput[59]), .A2(PermutationOutput[58]), .ZN(\Red_SubCellInst_LFInst_14_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_14_LFInst_1_U4  ( .A1(PermutationOutput[58]), 
        .A2(\Red_SubCellInst_LFInst_14_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_1_U3  ( .A(PermutationOutput[56]), 
        .B(PermutationOutput[59]), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_14_LFInst_2_n18 ), .ZN(Red_Feedback[58]) );
  AND2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_2_n17 ), .A2(PermutationOutput[56]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U8  ( .A1(PermutationOutput[58]), 
        .A2(PermutationOutput[57]), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_14_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_14_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U6  ( .A1(PermutationOutput[59]), 
        .A2(\Red_SubCellInst_LFInst_14_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U5  ( .A(PermutationOutput[57]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U4  ( .A1(PermutationOutput[58]), .A2(\Red_SubCellInst_LFInst_14_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U3  ( .A(PermutationOutput[56]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_3_U6  ( .A(PermutationOutput[57]), 
        .B(\Red_SubCellInst_LFInst_14_LFInst_3_n8 ), .ZN(Red_Feedback[59]) );
  NOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_14_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_3_U4  ( .A1(PermutationOutput[58]), 
        .A2(PermutationOutput[59]), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_14_LFInst_3_U3  ( .A1(PermutationOutput[59]), 
        .A2(PermutationOutput[56]), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_15_LFInst_0_n13 ), .ZN(Red_Feedback[60]) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U9  ( .A1(PermutationOutput[60]), .A2(\Red_SubCellInst_LFInst_15_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_0_n11 ), .A2(PermutationOutput[62]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_15_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_15_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U6  ( .A1(PermutationOutput[63]), .A2(\Red_SubCellInst_LFInst_15_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U5  ( .A(PermutationOutput[61]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U4  ( .A1(PermutationOutput[62]), .A2(\Red_SubCellInst_LFInst_15_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U3  ( .A(PermutationOutput[60]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_15_LFInst_1_n14 ), .ZN(Red_Feedback[61]) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_1_n13 ), .A2(PermutationOutput[61]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_1_n12 ), .A2(PermutationOutput[60]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_1_U5  ( .A1(PermutationOutput[63]), .A2(PermutationOutput[62]), .ZN(\Red_SubCellInst_LFInst_15_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_15_LFInst_1_U4  ( .A1(PermutationOutput[62]), 
        .A2(\Red_SubCellInst_LFInst_15_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_1_U3  ( .A(PermutationOutput[60]), 
        .B(PermutationOutput[63]), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_15_LFInst_2_n18 ), .ZN(Red_Feedback[62]) );
  AND2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_2_n17 ), .A2(PermutationOutput[60]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U8  ( .A1(PermutationOutput[62]), 
        .A2(PermutationOutput[61]), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_15_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_15_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U6  ( .A1(PermutationOutput[63]), 
        .A2(\Red_SubCellInst_LFInst_15_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U5  ( .A(PermutationOutput[61]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U4  ( .A1(PermutationOutput[62]), .A2(\Red_SubCellInst_LFInst_15_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U3  ( .A(PermutationOutput[60]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_3_U6  ( .A(PermutationOutput[61]), 
        .B(\Red_SubCellInst_LFInst_15_LFInst_3_n8 ), .ZN(Red_Feedback[63]) );
  NOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_15_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_3_U4  ( .A1(PermutationOutput[62]), 
        .A2(PermutationOutput[63]), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_15_LFInst_3_U3  ( .A1(PermutationOutput[63]), 
        .A2(PermutationOutput[60]), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_3_n7 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_0_LFInst_0_n2 ), .B(Key[2]), .ZN(Red_K0[0]) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_0_U3  ( .A(Key[3]), .B(Key[1]), .ZN(
        \Red_K0Inst_LFInst_0_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_0_LFInst_1_n2 ), .B(Key[2]), .ZN(Red_K0[1]) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_1_U3  ( .A(Key[3]), .B(Key[0]), .ZN(
        \Red_K0Inst_LFInst_0_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_0_LFInst_2_n2 ), .B(Key[1]), .ZN(Red_K0[2]) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_2_U3  ( .A(Key[3]), .B(Key[0]), .ZN(
        \Red_K0Inst_LFInst_0_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_0_LFInst_3_n2 ), .B(Key[1]), .ZN(Red_K0[3]) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_3_U3  ( .A(Key[2]), .B(Key[0]), .ZN(
        \Red_K0Inst_LFInst_0_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_1_LFInst_0_n2 ), .B(Key[6]), .ZN(Red_K0[4]) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_0_U3  ( .A(Key[7]), .B(Key[5]), .ZN(
        \Red_K0Inst_LFInst_1_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_1_LFInst_1_n2 ), .B(Key[6]), .ZN(Red_K0[5]) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_1_U3  ( .A(Key[7]), .B(Key[4]), .ZN(
        \Red_K0Inst_LFInst_1_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_1_LFInst_2_n2 ), .B(Key[5]), .ZN(Red_K0[6]) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_2_U3  ( .A(Key[7]), .B(Key[4]), .ZN(
        \Red_K0Inst_LFInst_1_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_1_LFInst_3_n2 ), .B(Key[5]), .ZN(Red_K0[7]) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_3_U3  ( .A(Key[6]), .B(Key[4]), .ZN(
        \Red_K0Inst_LFInst_1_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_2_LFInst_0_n2 ), .B(Key[10]), .ZN(Red_K0[8]) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_0_U3  ( .A(Key[11]), .B(Key[9]), .ZN(
        \Red_K0Inst_LFInst_2_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_2_LFInst_1_n2 ), .B(Key[10]), .ZN(Red_K0[9]) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_1_U3  ( .A(Key[11]), .B(Key[8]), .ZN(
        \Red_K0Inst_LFInst_2_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_2_LFInst_2_n2 ), .B(Key[9]), .ZN(Red_K0[10]) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_2_U3  ( .A(Key[11]), .B(Key[8]), .ZN(
        \Red_K0Inst_LFInst_2_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_2_LFInst_3_n2 ), .B(Key[9]), .ZN(Red_K0[11]) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_3_U3  ( .A(Key[10]), .B(Key[8]), .ZN(
        \Red_K0Inst_LFInst_2_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_3_LFInst_0_n2 ), .B(Key[14]), .ZN(Red_K0[12]) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_0_U3  ( .A(Key[15]), .B(Key[13]), .ZN(
        \Red_K0Inst_LFInst_3_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_3_LFInst_1_n2 ), .B(Key[14]), .ZN(Red_K0[13]) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_1_U3  ( .A(Key[15]), .B(Key[12]), .ZN(
        \Red_K0Inst_LFInst_3_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_3_LFInst_2_n2 ), .B(Key[13]), .ZN(Red_K0[14]) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_2_U3  ( .A(Key[15]), .B(Key[12]), .ZN(
        \Red_K0Inst_LFInst_3_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_3_LFInst_3_n2 ), .B(Key[13]), .ZN(Red_K0[15]) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_3_U3  ( .A(Key[14]), .B(Key[12]), .ZN(
        \Red_K0Inst_LFInst_3_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_4_LFInst_0_n2 ), .B(Key[18]), .ZN(Red_K0[16]) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_0_U3  ( .A(Key[19]), .B(Key[17]), .ZN(
        \Red_K0Inst_LFInst_4_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_4_LFInst_1_n2 ), .B(Key[18]), .ZN(Red_K0[17]) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_1_U3  ( .A(Key[19]), .B(Key[16]), .ZN(
        \Red_K0Inst_LFInst_4_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_4_LFInst_2_n2 ), .B(Key[17]), .ZN(Red_K0[18]) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_2_U3  ( .A(Key[19]), .B(Key[16]), .ZN(
        \Red_K0Inst_LFInst_4_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_4_LFInst_3_n2 ), .B(Key[17]), .ZN(Red_K0[19]) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_3_U3  ( .A(Key[18]), .B(Key[16]), .ZN(
        \Red_K0Inst_LFInst_4_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_5_LFInst_0_n2 ), .B(Key[22]), .ZN(Red_K0[20]) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_0_U3  ( .A(Key[23]), .B(Key[21]), .ZN(
        \Red_K0Inst_LFInst_5_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_5_LFInst_1_n2 ), .B(Key[22]), .ZN(Red_K0[21]) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_1_U3  ( .A(Key[23]), .B(Key[20]), .ZN(
        \Red_K0Inst_LFInst_5_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_5_LFInst_2_n2 ), .B(Key[21]), .ZN(Red_K0[22]) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_2_U3  ( .A(Key[23]), .B(Key[20]), .ZN(
        \Red_K0Inst_LFInst_5_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_5_LFInst_3_n2 ), .B(Key[21]), .ZN(Red_K0[23]) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_3_U3  ( .A(Key[22]), .B(Key[20]), .ZN(
        \Red_K0Inst_LFInst_5_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_6_LFInst_0_n2 ), .B(Key[26]), .ZN(Red_K0[24]) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_0_U3  ( .A(Key[27]), .B(Key[25]), .ZN(
        \Red_K0Inst_LFInst_6_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_6_LFInst_1_n2 ), .B(Key[26]), .ZN(Red_K0[25]) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_1_U3  ( .A(Key[27]), .B(Key[24]), .ZN(
        \Red_K0Inst_LFInst_6_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_6_LFInst_2_n2 ), .B(Key[25]), .ZN(Red_K0[26]) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_2_U3  ( .A(Key[27]), .B(Key[24]), .ZN(
        \Red_K0Inst_LFInst_6_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_6_LFInst_3_n2 ), .B(Key[25]), .ZN(Red_K0[27]) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_3_U3  ( .A(Key[26]), .B(Key[24]), .ZN(
        \Red_K0Inst_LFInst_6_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_7_LFInst_0_n2 ), .B(Key[30]), .ZN(Red_K0[28]) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_0_U3  ( .A(Key[31]), .B(Key[29]), .ZN(
        \Red_K0Inst_LFInst_7_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_7_LFInst_1_n2 ), .B(Key[30]), .ZN(Red_K0[29]) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_1_U3  ( .A(Key[31]), .B(Key[28]), .ZN(
        \Red_K0Inst_LFInst_7_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_7_LFInst_2_n2 ), .B(Key[29]), .ZN(Red_K0[30]) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_2_U3  ( .A(Key[31]), .B(Key[28]), .ZN(
        \Red_K0Inst_LFInst_7_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_7_LFInst_3_n2 ), .B(Key[29]), .ZN(Red_K0[31]) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_3_U3  ( .A(Key[30]), .B(Key[28]), .ZN(
        \Red_K0Inst_LFInst_7_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_8_LFInst_0_n2 ), .B(Key[34]), .ZN(Red_K0[32]) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_0_U3  ( .A(Key[35]), .B(Key[33]), .ZN(
        \Red_K0Inst_LFInst_8_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_8_LFInst_1_n2 ), .B(Key[34]), .ZN(Red_K0[33]) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_1_U3  ( .A(Key[35]), .B(Key[32]), .ZN(
        \Red_K0Inst_LFInst_8_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_8_LFInst_2_n2 ), .B(Key[33]), .ZN(Red_K0[34]) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_2_U3  ( .A(Key[35]), .B(Key[32]), .ZN(
        \Red_K0Inst_LFInst_8_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_8_LFInst_3_n2 ), .B(Key[33]), .ZN(Red_K0[35]) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_3_U3  ( .A(Key[34]), .B(Key[32]), .ZN(
        \Red_K0Inst_LFInst_8_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_9_LFInst_0_n2 ), .B(Key[38]), .ZN(Red_K0[36]) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_0_U3  ( .A(Key[39]), .B(Key[37]), .ZN(
        \Red_K0Inst_LFInst_9_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_9_LFInst_1_n2 ), .B(Key[38]), .ZN(Red_K0[37]) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_1_U3  ( .A(Key[39]), .B(Key[36]), .ZN(
        \Red_K0Inst_LFInst_9_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_9_LFInst_2_n2 ), .B(Key[37]), .ZN(Red_K0[38]) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_2_U3  ( .A(Key[39]), .B(Key[36]), .ZN(
        \Red_K0Inst_LFInst_9_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_9_LFInst_3_n2 ), .B(Key[37]), .ZN(Red_K0[39]) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_3_U3  ( .A(Key[38]), .B(Key[36]), .ZN(
        \Red_K0Inst_LFInst_9_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_10_LFInst_0_n2 ), .B(Key[42]), .ZN(Red_K0[40]) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_0_U3  ( .A(Key[43]), .B(Key[41]), .ZN(
        \Red_K0Inst_LFInst_10_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_10_LFInst_1_n2 ), .B(Key[42]), .ZN(Red_K0[41]) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_1_U3  ( .A(Key[43]), .B(Key[40]), .ZN(
        \Red_K0Inst_LFInst_10_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_10_LFInst_2_n2 ), .B(Key[41]), .ZN(Red_K0[42]) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_2_U3  ( .A(Key[43]), .B(Key[40]), .ZN(
        \Red_K0Inst_LFInst_10_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_10_LFInst_3_n2 ), .B(Key[41]), .ZN(Red_K0[43]) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_3_U3  ( .A(Key[42]), .B(Key[40]), .ZN(
        \Red_K0Inst_LFInst_10_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_11_LFInst_0_n2 ), .B(Key[46]), .ZN(Red_K0[44]) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_0_U3  ( .A(Key[47]), .B(Key[45]), .ZN(
        \Red_K0Inst_LFInst_11_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_11_LFInst_1_n2 ), .B(Key[46]), .ZN(Red_K0[45]) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_1_U3  ( .A(Key[47]), .B(Key[44]), .ZN(
        \Red_K0Inst_LFInst_11_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_11_LFInst_2_n2 ), .B(Key[45]), .ZN(Red_K0[46]) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_2_U3  ( .A(Key[47]), .B(Key[44]), .ZN(
        \Red_K0Inst_LFInst_11_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_11_LFInst_3_n2 ), .B(Key[45]), .ZN(Red_K0[47]) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_3_U3  ( .A(Key[46]), .B(Key[44]), .ZN(
        \Red_K0Inst_LFInst_11_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_12_LFInst_0_n2 ), .B(Key[50]), .ZN(Red_K0[48]) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_0_U3  ( .A(Key[51]), .B(Key[49]), .ZN(
        \Red_K0Inst_LFInst_12_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_12_LFInst_1_n2 ), .B(Key[50]), .ZN(Red_K0[49]) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_1_U3  ( .A(Key[51]), .B(Key[48]), .ZN(
        \Red_K0Inst_LFInst_12_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_12_LFInst_2_n2 ), .B(Key[49]), .ZN(Red_K0[50]) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_2_U3  ( .A(Key[51]), .B(Key[48]), .ZN(
        \Red_K0Inst_LFInst_12_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_12_LFInst_3_n2 ), .B(Key[49]), .ZN(Red_K0[51]) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_3_U3  ( .A(Key[50]), .B(Key[48]), .ZN(
        \Red_K0Inst_LFInst_12_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_13_LFInst_0_n2 ), .B(Key[54]), .ZN(Red_K0[52]) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_0_U3  ( .A(Key[55]), .B(Key[53]), .ZN(
        \Red_K0Inst_LFInst_13_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_13_LFInst_1_n2 ), .B(Key[54]), .ZN(Red_K0[53]) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_1_U3  ( .A(Key[55]), .B(Key[52]), .ZN(
        \Red_K0Inst_LFInst_13_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_13_LFInst_2_n2 ), .B(Key[53]), .ZN(Red_K0[54]) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_2_U3  ( .A(Key[55]), .B(Key[52]), .ZN(
        \Red_K0Inst_LFInst_13_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_13_LFInst_3_n2 ), .B(Key[53]), .ZN(Red_K0[55]) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_3_U3  ( .A(Key[54]), .B(Key[52]), .ZN(
        \Red_K0Inst_LFInst_13_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_14_LFInst_0_n2 ), .B(Key[58]), .ZN(Red_K0[56]) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_0_U3  ( .A(Key[59]), .B(Key[57]), .ZN(
        \Red_K0Inst_LFInst_14_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_14_LFInst_1_n2 ), .B(Key[58]), .ZN(Red_K0[57]) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_1_U3  ( .A(Key[59]), .B(Key[56]), .ZN(
        \Red_K0Inst_LFInst_14_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_14_LFInst_2_n2 ), .B(Key[57]), .ZN(Red_K0[58]) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_2_U3  ( .A(Key[59]), .B(Key[56]), .ZN(
        \Red_K0Inst_LFInst_14_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_14_LFInst_3_n2 ), .B(Key[57]), .ZN(Red_K0[59]) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_3_U3  ( .A(Key[58]), .B(Key[56]), .ZN(
        \Red_K0Inst_LFInst_14_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_15_LFInst_0_n2 ), .B(Key[62]), .ZN(Red_K0[60]) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_0_U3  ( .A(Key[63]), .B(Key[61]), .ZN(
        \Red_K0Inst_LFInst_15_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_15_LFInst_1_n2 ), .B(Key[62]), .ZN(Red_K0[61]) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_1_U3  ( .A(Key[63]), .B(Key[60]), .ZN(
        \Red_K0Inst_LFInst_15_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_15_LFInst_2_n2 ), .B(Key[61]), .ZN(Red_K0[62]) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_2_U3  ( .A(Key[63]), .B(Key[60]), .ZN(
        \Red_K0Inst_LFInst_15_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_15_LFInst_3_n2 ), .B(Key[61]), .ZN(Red_K0[63]) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_3_U3  ( .A(Key[62]), .B(Key[60]), .ZN(
        \Red_K0Inst_LFInst_15_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_0_LFInst_0_n2 ), .B(AddRoundKeyOutput[2]), 
        .ZN(Red_SignaltoCheck[0]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_0_U3  ( .A(AddRoundKeyOutput[3]), 
        .B(AddRoundKeyOutput[1]), .ZN(\Red_ToCheckInst_LFInst_0_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_0_LFInst_1_n2 ), .B(AddRoundKeyOutput[2]), 
        .ZN(Red_SignaltoCheck[1]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_1_U3  ( .A(AddRoundKeyOutput[3]), 
        .B(AddRoundKeyOutput[0]), .ZN(\Red_ToCheckInst_LFInst_0_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_0_LFInst_2_n2 ), .B(AddRoundKeyOutput[1]), 
        .ZN(Red_SignaltoCheck[2]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_2_U3  ( .A(AddRoundKeyOutput[3]), 
        .B(AddRoundKeyOutput[0]), .ZN(\Red_ToCheckInst_LFInst_0_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_0_LFInst_3_n2 ), .B(AddRoundKeyOutput[1]), 
        .ZN(Red_SignaltoCheck[3]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_3_U3  ( .A(AddRoundKeyOutput[2]), 
        .B(AddRoundKeyOutput[0]), .ZN(\Red_ToCheckInst_LFInst_0_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_1_LFInst_0_n2 ), .B(AddRoundKeyOutput[6]), 
        .ZN(Red_SignaltoCheck[4]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_0_U3  ( .A(AddRoundKeyOutput[7]), 
        .B(AddRoundKeyOutput[5]), .ZN(\Red_ToCheckInst_LFInst_1_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_1_LFInst_1_n2 ), .B(AddRoundKeyOutput[6]), 
        .ZN(Red_SignaltoCheck[5]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_1_U3  ( .A(AddRoundKeyOutput[7]), 
        .B(AddRoundKeyOutput[4]), .ZN(\Red_ToCheckInst_LFInst_1_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_1_LFInst_2_n2 ), .B(AddRoundKeyOutput[5]), 
        .ZN(Red_SignaltoCheck[6]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_2_U3  ( .A(AddRoundKeyOutput[7]), 
        .B(AddRoundKeyOutput[4]), .ZN(\Red_ToCheckInst_LFInst_1_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_1_LFInst_3_n2 ), .B(AddRoundKeyOutput[5]), 
        .ZN(Red_SignaltoCheck[7]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_3_U3  ( .A(AddRoundKeyOutput[6]), 
        .B(AddRoundKeyOutput[4]), .ZN(\Red_ToCheckInst_LFInst_1_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_2_LFInst_0_n2 ), .B(AddRoundKeyOutput[10]), 
        .ZN(Red_SignaltoCheck[8]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_0_U3  ( .A(AddRoundKeyOutput[11]), 
        .B(AddRoundKeyOutput[9]), .ZN(\Red_ToCheckInst_LFInst_2_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_2_LFInst_1_n2 ), .B(AddRoundKeyOutput[10]), 
        .ZN(Red_SignaltoCheck[9]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_1_U3  ( .A(AddRoundKeyOutput[11]), 
        .B(AddRoundKeyOutput[8]), .ZN(\Red_ToCheckInst_LFInst_2_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_2_LFInst_2_n2 ), .B(AddRoundKeyOutput[9]), 
        .ZN(Red_SignaltoCheck[10]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_2_U3  ( .A(AddRoundKeyOutput[11]), 
        .B(AddRoundKeyOutput[8]), .ZN(\Red_ToCheckInst_LFInst_2_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_2_LFInst_3_n2 ), .B(AddRoundKeyOutput[9]), 
        .ZN(Red_SignaltoCheck[11]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_3_U3  ( .A(AddRoundKeyOutput[10]), 
        .B(AddRoundKeyOutput[8]), .ZN(\Red_ToCheckInst_LFInst_2_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_3_LFInst_0_n2 ), .B(AddRoundKeyOutput[14]), 
        .ZN(Red_SignaltoCheck[12]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_0_U3  ( .A(AddRoundKeyOutput[15]), 
        .B(AddRoundKeyOutput[13]), .ZN(\Red_ToCheckInst_LFInst_3_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_3_LFInst_1_n2 ), .B(AddRoundKeyOutput[14]), 
        .ZN(Red_SignaltoCheck[13]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_1_U3  ( .A(AddRoundKeyOutput[15]), 
        .B(AddRoundKeyOutput[12]), .ZN(\Red_ToCheckInst_LFInst_3_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_3_LFInst_2_n2 ), .B(AddRoundKeyOutput[13]), 
        .ZN(Red_SignaltoCheck[14]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_2_U3  ( .A(AddRoundKeyOutput[15]), 
        .B(AddRoundKeyOutput[12]), .ZN(\Red_ToCheckInst_LFInst_3_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_3_LFInst_3_n2 ), .B(AddRoundKeyOutput[13]), 
        .ZN(Red_SignaltoCheck[15]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_3_U3  ( .A(AddRoundKeyOutput[14]), 
        .B(AddRoundKeyOutput[12]), .ZN(\Red_ToCheckInst_LFInst_3_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_4_LFInst_0_n2 ), .B(AddRoundKeyOutput[18]), 
        .ZN(Red_SignaltoCheck[16]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_0_U3  ( .A(AddRoundKeyOutput[19]), 
        .B(AddRoundKeyOutput[17]), .ZN(\Red_ToCheckInst_LFInst_4_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_4_LFInst_1_n2 ), .B(AddRoundKeyOutput[18]), 
        .ZN(Red_SignaltoCheck[17]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_1_U3  ( .A(AddRoundKeyOutput[19]), 
        .B(AddRoundKeyOutput[16]), .ZN(\Red_ToCheckInst_LFInst_4_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_4_LFInst_2_n2 ), .B(AddRoundKeyOutput[17]), 
        .ZN(Red_SignaltoCheck[18]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_2_U3  ( .A(AddRoundKeyOutput[19]), 
        .B(AddRoundKeyOutput[16]), .ZN(\Red_ToCheckInst_LFInst_4_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_4_LFInst_3_n2 ), .B(AddRoundKeyOutput[17]), 
        .ZN(Red_SignaltoCheck[19]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_3_U3  ( .A(AddRoundKeyOutput[18]), 
        .B(AddRoundKeyOutput[16]), .ZN(\Red_ToCheckInst_LFInst_4_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_5_LFInst_0_n2 ), .B(AddRoundKeyOutput[22]), 
        .ZN(Red_SignaltoCheck[20]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_0_U3  ( .A(AddRoundKeyOutput[23]), 
        .B(AddRoundKeyOutput[21]), .ZN(\Red_ToCheckInst_LFInst_5_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_5_LFInst_1_n2 ), .B(AddRoundKeyOutput[22]), 
        .ZN(Red_SignaltoCheck[21]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_1_U3  ( .A(AddRoundKeyOutput[23]), 
        .B(AddRoundKeyOutput[20]), .ZN(\Red_ToCheckInst_LFInst_5_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_5_LFInst_2_n2 ), .B(AddRoundKeyOutput[21]), 
        .ZN(Red_SignaltoCheck[22]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_2_U3  ( .A(AddRoundKeyOutput[23]), 
        .B(AddRoundKeyOutput[20]), .ZN(\Red_ToCheckInst_LFInst_5_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_5_LFInst_3_n2 ), .B(AddRoundKeyOutput[21]), 
        .ZN(Red_SignaltoCheck[23]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_3_U3  ( .A(AddRoundKeyOutput[22]), 
        .B(AddRoundKeyOutput[20]), .ZN(\Red_ToCheckInst_LFInst_5_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_6_LFInst_0_n2 ), .B(AddRoundKeyOutput[26]), 
        .ZN(Red_SignaltoCheck[24]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_0_U3  ( .A(AddRoundKeyOutput[27]), 
        .B(AddRoundKeyOutput[25]), .ZN(\Red_ToCheckInst_LFInst_6_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_6_LFInst_1_n2 ), .B(AddRoundKeyOutput[26]), 
        .ZN(Red_SignaltoCheck[25]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_1_U3  ( .A(AddRoundKeyOutput[27]), 
        .B(AddRoundKeyOutput[24]), .ZN(\Red_ToCheckInst_LFInst_6_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_6_LFInst_2_n2 ), .B(AddRoundKeyOutput[25]), 
        .ZN(Red_SignaltoCheck[26]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_2_U3  ( .A(AddRoundKeyOutput[27]), 
        .B(AddRoundKeyOutput[24]), .ZN(\Red_ToCheckInst_LFInst_6_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_6_LFInst_3_n2 ), .B(AddRoundKeyOutput[25]), 
        .ZN(Red_SignaltoCheck[27]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_3_U3  ( .A(AddRoundKeyOutput[26]), 
        .B(AddRoundKeyOutput[24]), .ZN(\Red_ToCheckInst_LFInst_6_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_7_LFInst_0_n2 ), .B(AddRoundKeyOutput[30]), 
        .ZN(Red_SignaltoCheck[28]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_0_U3  ( .A(AddRoundKeyOutput[31]), 
        .B(AddRoundKeyOutput[29]), .ZN(\Red_ToCheckInst_LFInst_7_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_7_LFInst_1_n2 ), .B(AddRoundKeyOutput[30]), 
        .ZN(Red_SignaltoCheck[29]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_1_U3  ( .A(AddRoundKeyOutput[31]), 
        .B(AddRoundKeyOutput[28]), .ZN(\Red_ToCheckInst_LFInst_7_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_7_LFInst_2_n2 ), .B(AddRoundKeyOutput[29]), 
        .ZN(Red_SignaltoCheck[30]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_2_U3  ( .A(AddRoundKeyOutput[31]), 
        .B(AddRoundKeyOutput[28]), .ZN(\Red_ToCheckInst_LFInst_7_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_7_LFInst_3_n2 ), .B(AddRoundKeyOutput[29]), 
        .ZN(Red_SignaltoCheck[31]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_3_U3  ( .A(AddRoundKeyOutput[30]), 
        .B(AddRoundKeyOutput[28]), .ZN(\Red_ToCheckInst_LFInst_7_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_8_LFInst_0_n2 ), .B(AddRoundKeyOutput[34]), 
        .ZN(Red_SignaltoCheck[32]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_0_U3  ( .A(AddRoundKeyOutput[35]), 
        .B(AddRoundKeyOutput[33]), .ZN(\Red_ToCheckInst_LFInst_8_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_8_LFInst_1_n2 ), .B(AddRoundKeyOutput[34]), 
        .ZN(Red_SignaltoCheck[33]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_1_U3  ( .A(AddRoundKeyOutput[35]), 
        .B(AddRoundKeyOutput[32]), .ZN(\Red_ToCheckInst_LFInst_8_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_8_LFInst_2_n2 ), .B(AddRoundKeyOutput[33]), 
        .ZN(Red_SignaltoCheck[34]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_2_U3  ( .A(AddRoundKeyOutput[35]), 
        .B(AddRoundKeyOutput[32]), .ZN(\Red_ToCheckInst_LFInst_8_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_8_LFInst_3_n2 ), .B(AddRoundKeyOutput[33]), 
        .ZN(Red_SignaltoCheck[35]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_3_U3  ( .A(AddRoundKeyOutput[34]), 
        .B(AddRoundKeyOutput[32]), .ZN(\Red_ToCheckInst_LFInst_8_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_9_LFInst_0_n2 ), .B(AddRoundKeyOutput[38]), 
        .ZN(Red_SignaltoCheck[36]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_0_U3  ( .A(AddRoundKeyOutput[39]), 
        .B(AddRoundKeyOutput[37]), .ZN(\Red_ToCheckInst_LFInst_9_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_9_LFInst_1_n2 ), .B(AddRoundKeyOutput[38]), 
        .ZN(Red_SignaltoCheck[37]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_1_U3  ( .A(AddRoundKeyOutput[39]), 
        .B(AddRoundKeyOutput[36]), .ZN(\Red_ToCheckInst_LFInst_9_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_9_LFInst_2_n2 ), .B(AddRoundKeyOutput[37]), 
        .ZN(Red_SignaltoCheck[38]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_2_U3  ( .A(AddRoundKeyOutput[39]), 
        .B(AddRoundKeyOutput[36]), .ZN(\Red_ToCheckInst_LFInst_9_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_9_LFInst_3_n2 ), .B(AddRoundKeyOutput[37]), 
        .ZN(Red_SignaltoCheck[39]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_3_U3  ( .A(AddRoundKeyOutput[38]), 
        .B(AddRoundKeyOutput[36]), .ZN(\Red_ToCheckInst_LFInst_9_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_10_LFInst_0_n2 ), .B(AddRoundKeyOutput[42]), 
        .ZN(Red_SignaltoCheck[40]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_0_U3  ( .A(AddRoundKeyOutput[43]), 
        .B(AddRoundKeyOutput[41]), .ZN(\Red_ToCheckInst_LFInst_10_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_10_LFInst_1_n2 ), .B(AddRoundKeyOutput[42]), 
        .ZN(Red_SignaltoCheck[41]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_1_U3  ( .A(AddRoundKeyOutput[43]), 
        .B(AddRoundKeyOutput[40]), .ZN(\Red_ToCheckInst_LFInst_10_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_10_LFInst_2_n2 ), .B(AddRoundKeyOutput[41]), 
        .ZN(Red_SignaltoCheck[42]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_2_U3  ( .A(AddRoundKeyOutput[43]), 
        .B(AddRoundKeyOutput[40]), .ZN(\Red_ToCheckInst_LFInst_10_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_10_LFInst_3_n2 ), .B(AddRoundKeyOutput[41]), 
        .ZN(Red_SignaltoCheck[43]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_3_U3  ( .A(AddRoundKeyOutput[42]), 
        .B(AddRoundKeyOutput[40]), .ZN(\Red_ToCheckInst_LFInst_10_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_11_LFInst_0_n2 ), .B(AddRoundKeyOutput[46]), 
        .ZN(Red_SignaltoCheck[44]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_0_U3  ( .A(AddRoundKeyOutput[47]), 
        .B(AddRoundKeyOutput[45]), .ZN(\Red_ToCheckInst_LFInst_11_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_11_LFInst_1_n2 ), .B(AddRoundKeyOutput[46]), 
        .ZN(Red_SignaltoCheck[45]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_1_U3  ( .A(AddRoundKeyOutput[47]), 
        .B(AddRoundKeyOutput[44]), .ZN(\Red_ToCheckInst_LFInst_11_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_11_LFInst_2_n2 ), .B(AddRoundKeyOutput[45]), 
        .ZN(Red_SignaltoCheck[46]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_2_U3  ( .A(AddRoundKeyOutput[47]), 
        .B(AddRoundKeyOutput[44]), .ZN(\Red_ToCheckInst_LFInst_11_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_11_LFInst_3_n2 ), .B(AddRoundKeyOutput[45]), 
        .ZN(Red_SignaltoCheck[47]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_3_U3  ( .A(AddRoundKeyOutput[46]), 
        .B(AddRoundKeyOutput[44]), .ZN(\Red_ToCheckInst_LFInst_11_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_12_LFInst_0_n2 ), .B(AddRoundKeyOutput[50]), 
        .ZN(Red_SignaltoCheck[48]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_0_U3  ( .A(AddRoundKeyOutput[51]), 
        .B(AddRoundKeyOutput[49]), .ZN(\Red_ToCheckInst_LFInst_12_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_12_LFInst_1_n2 ), .B(AddRoundKeyOutput[50]), 
        .ZN(Red_SignaltoCheck[49]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_1_U3  ( .A(AddRoundKeyOutput[51]), 
        .B(AddRoundKeyOutput[48]), .ZN(\Red_ToCheckInst_LFInst_12_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_12_LFInst_2_n2 ), .B(AddRoundKeyOutput[49]), 
        .ZN(Red_SignaltoCheck[50]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_2_U3  ( .A(AddRoundKeyOutput[51]), 
        .B(AddRoundKeyOutput[48]), .ZN(\Red_ToCheckInst_LFInst_12_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_12_LFInst_3_n2 ), .B(AddRoundKeyOutput[49]), 
        .ZN(Red_SignaltoCheck[51]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_3_U3  ( .A(AddRoundKeyOutput[50]), 
        .B(AddRoundKeyOutput[48]), .ZN(\Red_ToCheckInst_LFInst_12_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_13_LFInst_0_n2 ), .B(AddRoundKeyOutput[54]), 
        .ZN(Red_SignaltoCheck[52]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_0_U3  ( .A(AddRoundKeyOutput[55]), 
        .B(AddRoundKeyOutput[53]), .ZN(\Red_ToCheckInst_LFInst_13_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_13_LFInst_1_n2 ), .B(AddRoundKeyOutput[54]), 
        .ZN(Red_SignaltoCheck[53]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_1_U3  ( .A(AddRoundKeyOutput[55]), 
        .B(AddRoundKeyOutput[52]), .ZN(\Red_ToCheckInst_LFInst_13_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_13_LFInst_2_n2 ), .B(AddRoundKeyOutput[53]), 
        .ZN(Red_SignaltoCheck[54]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_2_U3  ( .A(AddRoundKeyOutput[55]), 
        .B(AddRoundKeyOutput[52]), .ZN(\Red_ToCheckInst_LFInst_13_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_13_LFInst_3_n2 ), .B(AddRoundKeyOutput[53]), 
        .ZN(Red_SignaltoCheck[55]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_3_U3  ( .A(AddRoundKeyOutput[54]), 
        .B(AddRoundKeyOutput[52]), .ZN(\Red_ToCheckInst_LFInst_13_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_14_LFInst_0_n2 ), .B(AddRoundKeyOutput[58]), 
        .ZN(Red_SignaltoCheck[56]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_0_U3  ( .A(AddRoundKeyOutput[59]), 
        .B(AddRoundKeyOutput[57]), .ZN(\Red_ToCheckInst_LFInst_14_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_14_LFInst_1_n2 ), .B(AddRoundKeyOutput[58]), 
        .ZN(Red_SignaltoCheck[57]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_1_U3  ( .A(AddRoundKeyOutput[59]), 
        .B(AddRoundKeyOutput[56]), .ZN(\Red_ToCheckInst_LFInst_14_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_14_LFInst_2_n2 ), .B(AddRoundKeyOutput[57]), 
        .ZN(Red_SignaltoCheck[58]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_2_U3  ( .A(AddRoundKeyOutput[59]), 
        .B(AddRoundKeyOutput[56]), .ZN(\Red_ToCheckInst_LFInst_14_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_14_LFInst_3_n2 ), .B(AddRoundKeyOutput[57]), 
        .ZN(Red_SignaltoCheck[59]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_3_U3  ( .A(AddRoundKeyOutput[58]), 
        .B(AddRoundKeyOutput[56]), .ZN(\Red_ToCheckInst_LFInst_14_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_15_LFInst_0_n2 ), .B(AddRoundKeyOutput[62]), 
        .ZN(Red_SignaltoCheck[60]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_0_U3  ( .A(AddRoundKeyOutput[63]), 
        .B(AddRoundKeyOutput[61]), .ZN(\Red_ToCheckInst_LFInst_15_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_15_LFInst_1_n2 ), .B(AddRoundKeyOutput[62]), 
        .ZN(Red_SignaltoCheck[61]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_1_U3  ( .A(AddRoundKeyOutput[63]), 
        .B(AddRoundKeyOutput[60]), .ZN(\Red_ToCheckInst_LFInst_15_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_15_LFInst_2_n2 ), .B(AddRoundKeyOutput[61]), 
        .ZN(Red_SignaltoCheck[62]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_2_U3  ( .A(AddRoundKeyOutput[63]), 
        .B(AddRoundKeyOutput[60]), .ZN(\Red_ToCheckInst_LFInst_15_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_15_LFInst_3_n2 ), .B(AddRoundKeyOutput[61]), 
        .ZN(Red_SignaltoCheck[63]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_3_U3  ( .A(AddRoundKeyOutput[62]), 
        .B(AddRoundKeyOutput[60]), .ZN(\Red_ToCheckInst_LFInst_15_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_16_LFInst_0_n2 ), .B(Output[2]), .ZN(
        Red_SignaltoCheck[64]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_0_U3  ( .A(Output[3]), .B(
        Output[1]), .ZN(\Red_ToCheckInst_LFInst_16_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_16_LFInst_1_n2 ), .B(Output[2]), .ZN(
        Red_SignaltoCheck[65]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_1_U3  ( .A(Output[3]), .B(
        Output[0]), .ZN(\Red_ToCheckInst_LFInst_16_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_16_LFInst_2_n2 ), .B(Output[1]), .ZN(
        Red_SignaltoCheck[66]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_2_U3  ( .A(Output[3]), .B(
        Output[0]), .ZN(\Red_ToCheckInst_LFInst_16_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_16_LFInst_3_n2 ), .B(Output[1]), .ZN(
        Red_SignaltoCheck[67]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_3_U3  ( .A(Output[2]), .B(
        Output[0]), .ZN(\Red_ToCheckInst_LFInst_16_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_17_LFInst_0_n2 ), .B(Output[6]), .ZN(
        Red_SignaltoCheck[68]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_0_U3  ( .A(Output[7]), .B(
        Output[5]), .ZN(\Red_ToCheckInst_LFInst_17_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_17_LFInst_1_n2 ), .B(Output[6]), .ZN(
        Red_SignaltoCheck[69]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_1_U3  ( .A(Output[7]), .B(
        Output[4]), .ZN(\Red_ToCheckInst_LFInst_17_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_17_LFInst_2_n2 ), .B(Output[5]), .ZN(
        Red_SignaltoCheck[70]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_2_U3  ( .A(Output[7]), .B(
        Output[4]), .ZN(\Red_ToCheckInst_LFInst_17_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_17_LFInst_3_n2 ), .B(Output[5]), .ZN(
        Red_SignaltoCheck[71]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_3_U3  ( .A(Output[6]), .B(
        Output[4]), .ZN(\Red_ToCheckInst_LFInst_17_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_18_LFInst_0_n2 ), .B(Output[10]), .ZN(
        Red_SignaltoCheck[72]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_0_U3  ( .A(Output[11]), .B(
        Output[9]), .ZN(\Red_ToCheckInst_LFInst_18_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_18_LFInst_1_n2 ), .B(Output[10]), .ZN(
        Red_SignaltoCheck[73]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_1_U3  ( .A(Output[11]), .B(
        Output[8]), .ZN(\Red_ToCheckInst_LFInst_18_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_18_LFInst_2_n2 ), .B(Output[9]), .ZN(
        Red_SignaltoCheck[74]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_2_U3  ( .A(Output[11]), .B(
        Output[8]), .ZN(\Red_ToCheckInst_LFInst_18_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_18_LFInst_3_n2 ), .B(Output[9]), .ZN(
        Red_SignaltoCheck[75]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_3_U3  ( .A(Output[10]), .B(
        Output[8]), .ZN(\Red_ToCheckInst_LFInst_18_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_19_LFInst_0_n2 ), .B(Output[14]), .ZN(
        Red_SignaltoCheck[76]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_0_U3  ( .A(Output[15]), .B(
        Output[13]), .ZN(\Red_ToCheckInst_LFInst_19_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_19_LFInst_1_n2 ), .B(Output[14]), .ZN(
        Red_SignaltoCheck[77]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_1_U3  ( .A(Output[15]), .B(
        Output[12]), .ZN(\Red_ToCheckInst_LFInst_19_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_19_LFInst_2_n2 ), .B(Output[13]), .ZN(
        Red_SignaltoCheck[78]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_2_U3  ( .A(Output[15]), .B(
        Output[12]), .ZN(\Red_ToCheckInst_LFInst_19_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_19_LFInst_3_n2 ), .B(Output[13]), .ZN(
        Red_SignaltoCheck[79]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_3_U3  ( .A(Output[14]), .B(
        Output[12]), .ZN(\Red_ToCheckInst_LFInst_19_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_20_LFInst_0_n2 ), .B(Output[18]), .ZN(
        Red_SignaltoCheck[80]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_0_U3  ( .A(Output[19]), .B(
        Output[17]), .ZN(\Red_ToCheckInst_LFInst_20_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_20_LFInst_1_n2 ), .B(Output[18]), .ZN(
        Red_SignaltoCheck[81]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_1_U3  ( .A(Output[19]), .B(
        Output[16]), .ZN(\Red_ToCheckInst_LFInst_20_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_20_LFInst_2_n2 ), .B(Output[17]), .ZN(
        Red_SignaltoCheck[82]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_2_U3  ( .A(Output[19]), .B(
        Output[16]), .ZN(\Red_ToCheckInst_LFInst_20_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_20_LFInst_3_n2 ), .B(Output[17]), .ZN(
        Red_SignaltoCheck[83]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_3_U3  ( .A(Output[18]), .B(
        Output[16]), .ZN(\Red_ToCheckInst_LFInst_20_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_21_LFInst_0_n2 ), .B(Output[22]), .ZN(
        Red_SignaltoCheck[84]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_0_U3  ( .A(Output[23]), .B(
        Output[21]), .ZN(\Red_ToCheckInst_LFInst_21_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_21_LFInst_1_n2 ), .B(Output[22]), .ZN(
        Red_SignaltoCheck[85]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_1_U3  ( .A(Output[23]), .B(
        Output[20]), .ZN(\Red_ToCheckInst_LFInst_21_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_21_LFInst_2_n2 ), .B(Output[21]), .ZN(
        Red_SignaltoCheck[86]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_2_U3  ( .A(Output[23]), .B(
        Output[20]), .ZN(\Red_ToCheckInst_LFInst_21_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_21_LFInst_3_n2 ), .B(Output[21]), .ZN(
        Red_SignaltoCheck[87]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_3_U3  ( .A(Output[22]), .B(
        Output[20]), .ZN(\Red_ToCheckInst_LFInst_21_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_22_LFInst_0_n2 ), .B(Output[26]), .ZN(
        Red_SignaltoCheck[88]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_0_U3  ( .A(Output[27]), .B(
        Output[25]), .ZN(\Red_ToCheckInst_LFInst_22_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_22_LFInst_1_n2 ), .B(Output[26]), .ZN(
        Red_SignaltoCheck[89]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_1_U3  ( .A(Output[27]), .B(
        Output[24]), .ZN(\Red_ToCheckInst_LFInst_22_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_22_LFInst_2_n2 ), .B(Output[25]), .ZN(
        Red_SignaltoCheck[90]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_2_U3  ( .A(Output[27]), .B(
        Output[24]), .ZN(\Red_ToCheckInst_LFInst_22_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_22_LFInst_3_n2 ), .B(Output[25]), .ZN(
        Red_SignaltoCheck[91]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_3_U3  ( .A(Output[26]), .B(
        Output[24]), .ZN(\Red_ToCheckInst_LFInst_22_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_23_LFInst_0_n2 ), .B(Output[30]), .ZN(
        Red_SignaltoCheck[92]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_0_U3  ( .A(Output[31]), .B(
        Output[29]), .ZN(\Red_ToCheckInst_LFInst_23_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_23_LFInst_1_n2 ), .B(Output[30]), .ZN(
        Red_SignaltoCheck[93]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_1_U3  ( .A(Output[31]), .B(
        Output[28]), .ZN(\Red_ToCheckInst_LFInst_23_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_23_LFInst_2_n2 ), .B(Output[29]), .ZN(
        Red_SignaltoCheck[94]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_2_U3  ( .A(Output[31]), .B(
        Output[28]), .ZN(\Red_ToCheckInst_LFInst_23_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_23_LFInst_3_n2 ), .B(Output[29]), .ZN(
        Red_SignaltoCheck[95]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_3_U3  ( .A(Output[30]), .B(
        Output[28]), .ZN(\Red_ToCheckInst_LFInst_23_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_24_LFInst_0_n2 ), .B(Output[34]), .ZN(
        Red_SignaltoCheck[96]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_0_U3  ( .A(Output[35]), .B(
        Output[33]), .ZN(\Red_ToCheckInst_LFInst_24_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_24_LFInst_1_n2 ), .B(Output[34]), .ZN(
        Red_SignaltoCheck[97]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_1_U3  ( .A(Output[35]), .B(
        Output[32]), .ZN(\Red_ToCheckInst_LFInst_24_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_24_LFInst_2_n2 ), .B(Output[33]), .ZN(
        Red_SignaltoCheck[98]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_2_U3  ( .A(Output[35]), .B(
        Output[32]), .ZN(\Red_ToCheckInst_LFInst_24_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_24_LFInst_3_n2 ), .B(Output[33]), .ZN(
        Red_SignaltoCheck[99]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_3_U3  ( .A(Output[34]), .B(
        Output[32]), .ZN(\Red_ToCheckInst_LFInst_24_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_25_LFInst_0_n2 ), .B(Output[38]), .ZN(
        Red_SignaltoCheck[100]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_0_U3  ( .A(Output[39]), .B(
        Output[37]), .ZN(\Red_ToCheckInst_LFInst_25_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_25_LFInst_1_n2 ), .B(Output[38]), .ZN(
        Red_SignaltoCheck[101]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_1_U3  ( .A(Output[39]), .B(
        Output[36]), .ZN(\Red_ToCheckInst_LFInst_25_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_25_LFInst_2_n2 ), .B(Output[37]), .ZN(
        Red_SignaltoCheck[102]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_2_U3  ( .A(Output[39]), .B(
        Output[36]), .ZN(\Red_ToCheckInst_LFInst_25_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_25_LFInst_3_n2 ), .B(Output[37]), .ZN(
        Red_SignaltoCheck[103]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_3_U3  ( .A(Output[38]), .B(
        Output[36]), .ZN(\Red_ToCheckInst_LFInst_25_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_26_LFInst_0_n2 ), .B(Output[42]), .ZN(
        Red_SignaltoCheck[104]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_0_U3  ( .A(Output[43]), .B(
        Output[41]), .ZN(\Red_ToCheckInst_LFInst_26_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_26_LFInst_1_n2 ), .B(Output[42]), .ZN(
        Red_SignaltoCheck[105]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_1_U3  ( .A(Output[43]), .B(
        Output[40]), .ZN(\Red_ToCheckInst_LFInst_26_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_26_LFInst_2_n2 ), .B(Output[41]), .ZN(
        Red_SignaltoCheck[106]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_2_U3  ( .A(Output[43]), .B(
        Output[40]), .ZN(\Red_ToCheckInst_LFInst_26_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_26_LFInst_3_n2 ), .B(Output[41]), .ZN(
        Red_SignaltoCheck[107]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_3_U3  ( .A(Output[42]), .B(
        Output[40]), .ZN(\Red_ToCheckInst_LFInst_26_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_27_LFInst_0_n2 ), .B(Output[46]), .ZN(
        Red_SignaltoCheck[108]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_0_U3  ( .A(Output[47]), .B(
        Output[45]), .ZN(\Red_ToCheckInst_LFInst_27_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_27_LFInst_1_n2 ), .B(Output[46]), .ZN(
        Red_SignaltoCheck[109]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_1_U3  ( .A(Output[47]), .B(
        Output[44]), .ZN(\Red_ToCheckInst_LFInst_27_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_27_LFInst_2_n2 ), .B(Output[45]), .ZN(
        Red_SignaltoCheck[110]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_2_U3  ( .A(Output[47]), .B(
        Output[44]), .ZN(\Red_ToCheckInst_LFInst_27_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_27_LFInst_3_n2 ), .B(Output[45]), .ZN(
        Red_SignaltoCheck[111]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_3_U3  ( .A(Output[46]), .B(
        Output[44]), .ZN(\Red_ToCheckInst_LFInst_27_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_28_LFInst_0_n2 ), .B(Output[50]), .ZN(
        Red_SignaltoCheck[112]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_0_U3  ( .A(Output[51]), .B(
        Output[49]), .ZN(\Red_ToCheckInst_LFInst_28_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_28_LFInst_1_n2 ), .B(Output[50]), .ZN(
        Red_SignaltoCheck[113]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_1_U3  ( .A(Output[51]), .B(
        Output[48]), .ZN(\Red_ToCheckInst_LFInst_28_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_28_LFInst_2_n2 ), .B(Output[49]), .ZN(
        Red_SignaltoCheck[114]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_2_U3  ( .A(Output[51]), .B(
        Output[48]), .ZN(\Red_ToCheckInst_LFInst_28_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_28_LFInst_3_n2 ), .B(Output[49]), .ZN(
        Red_SignaltoCheck[115]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_3_U3  ( .A(Output[50]), .B(
        Output[48]), .ZN(\Red_ToCheckInst_LFInst_28_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_29_LFInst_0_n2 ), .B(Output[54]), .ZN(
        Red_SignaltoCheck[116]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_0_U3  ( .A(Output[55]), .B(
        Output[53]), .ZN(\Red_ToCheckInst_LFInst_29_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_29_LFInst_1_n2 ), .B(Output[54]), .ZN(
        Red_SignaltoCheck[117]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_1_U3  ( .A(Output[55]), .B(
        Output[52]), .ZN(\Red_ToCheckInst_LFInst_29_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_29_LFInst_2_n2 ), .B(Output[53]), .ZN(
        Red_SignaltoCheck[118]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_2_U3  ( .A(Output[55]), .B(
        Output[52]), .ZN(\Red_ToCheckInst_LFInst_29_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_29_LFInst_3_n2 ), .B(Output[53]), .ZN(
        Red_SignaltoCheck[119]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_3_U3  ( .A(Output[54]), .B(
        Output[52]), .ZN(\Red_ToCheckInst_LFInst_29_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_30_LFInst_0_n2 ), .B(Output[58]), .ZN(
        Red_SignaltoCheck[120]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_0_U3  ( .A(Output[59]), .B(
        Output[57]), .ZN(\Red_ToCheckInst_LFInst_30_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_30_LFInst_1_n2 ), .B(Output[58]), .ZN(
        Red_SignaltoCheck[121]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_1_U3  ( .A(Output[59]), .B(
        Output[56]), .ZN(\Red_ToCheckInst_LFInst_30_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_30_LFInst_2_n2 ), .B(Output[57]), .ZN(
        Red_SignaltoCheck[122]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_2_U3  ( .A(Output[59]), .B(
        Output[56]), .ZN(\Red_ToCheckInst_LFInst_30_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_30_LFInst_3_n2 ), .B(Output[57]), .ZN(
        Red_SignaltoCheck[123]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_3_U3  ( .A(Output[58]), .B(
        Output[56]), .ZN(\Red_ToCheckInst_LFInst_30_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_31_LFInst_0_n2 ), .B(Output[62]), .ZN(
        Red_SignaltoCheck[124]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_0_U3  ( .A(Output[63]), .B(
        Output[61]), .ZN(\Red_ToCheckInst_LFInst_31_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_31_LFInst_1_n2 ), .B(Output[62]), .ZN(
        Red_SignaltoCheck[125]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_1_U3  ( .A(Output[63]), .B(
        Output[60]), .ZN(\Red_ToCheckInst_LFInst_31_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_31_LFInst_2_n2 ), .B(Output[61]), .ZN(
        Red_SignaltoCheck[126]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_2_U3  ( .A(Output[63]), .B(
        Output[60]), .ZN(\Red_ToCheckInst_LFInst_31_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_31_LFInst_3_n2 ), .B(Output[61]), .ZN(
        Red_SignaltoCheck[127]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_3_U3  ( .A(Output[62]), .B(
        Output[60]), .ZN(\Red_ToCheckInst_LFInst_31_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_32_LFInst_0_n2 ), .B(PermutationOutput[62]), 
        .ZN(Red_SignaltoCheck[128]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_0_U3  ( .A(PermutationOutput[63]), 
        .B(PermutationOutput[61]), .ZN(\Red_ToCheckInst_LFInst_32_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_32_LFInst_1_n2 ), .B(PermutationOutput[62]), 
        .ZN(Red_SignaltoCheck[129]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_1_U3  ( .A(PermutationOutput[63]), 
        .B(PermutationOutput[60]), .ZN(\Red_ToCheckInst_LFInst_32_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_32_LFInst_2_n2 ), .B(PermutationOutput[61]), 
        .ZN(Red_SignaltoCheck[130]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_2_U3  ( .A(PermutationOutput[63]), 
        .B(PermutationOutput[60]), .ZN(\Red_ToCheckInst_LFInst_32_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_32_LFInst_3_n2 ), .B(PermutationOutput[61]), 
        .ZN(Red_SignaltoCheck[131]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_3_U3  ( .A(PermutationOutput[62]), 
        .B(PermutationOutput[60]), .ZN(\Red_ToCheckInst_LFInst_32_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_33_LFInst_0_n2 ), .B(PermutationOutput[50]), 
        .ZN(Red_SignaltoCheck[132]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_0_U3  ( .A(PermutationOutput[51]), 
        .B(PermutationOutput[49]), .ZN(\Red_ToCheckInst_LFInst_33_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_33_LFInst_1_n2 ), .B(PermutationOutput[50]), 
        .ZN(Red_SignaltoCheck[133]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_1_U3  ( .A(PermutationOutput[51]), 
        .B(PermutationOutput[48]), .ZN(\Red_ToCheckInst_LFInst_33_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_33_LFInst_2_n2 ), .B(PermutationOutput[49]), 
        .ZN(Red_SignaltoCheck[134]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_2_U3  ( .A(PermutationOutput[51]), 
        .B(PermutationOutput[48]), .ZN(\Red_ToCheckInst_LFInst_33_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_33_LFInst_3_n2 ), .B(PermutationOutput[49]), 
        .ZN(Red_SignaltoCheck[135]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_3_U3  ( .A(PermutationOutput[50]), 
        .B(PermutationOutput[48]), .ZN(\Red_ToCheckInst_LFInst_33_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_34_LFInst_0_n2 ), .B(PermutationOutput[54]), 
        .ZN(Red_SignaltoCheck[136]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_0_U3  ( .A(PermutationOutput[55]), 
        .B(PermutationOutput[53]), .ZN(\Red_ToCheckInst_LFInst_34_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_34_LFInst_1_n2 ), .B(PermutationOutput[54]), 
        .ZN(Red_SignaltoCheck[137]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_1_U3  ( .A(PermutationOutput[55]), 
        .B(PermutationOutput[52]), .ZN(\Red_ToCheckInst_LFInst_34_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_34_LFInst_2_n2 ), .B(PermutationOutput[53]), 
        .ZN(Red_SignaltoCheck[138]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_2_U3  ( .A(PermutationOutput[55]), 
        .B(PermutationOutput[52]), .ZN(\Red_ToCheckInst_LFInst_34_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_34_LFInst_3_n2 ), .B(PermutationOutput[53]), 
        .ZN(Red_SignaltoCheck[139]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_3_U3  ( .A(PermutationOutput[54]), 
        .B(PermutationOutput[52]), .ZN(\Red_ToCheckInst_LFInst_34_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_35_LFInst_0_n2 ), .B(PermutationOutput[58]), 
        .ZN(Red_SignaltoCheck[140]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_0_U3  ( .A(PermutationOutput[59]), 
        .B(PermutationOutput[57]), .ZN(\Red_ToCheckInst_LFInst_35_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_35_LFInst_1_n2 ), .B(PermutationOutput[58]), 
        .ZN(Red_SignaltoCheck[141]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_1_U3  ( .A(PermutationOutput[59]), 
        .B(PermutationOutput[56]), .ZN(\Red_ToCheckInst_LFInst_35_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_35_LFInst_2_n2 ), .B(PermutationOutput[57]), 
        .ZN(Red_SignaltoCheck[142]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_2_U3  ( .A(PermutationOutput[59]), 
        .B(PermutationOutput[56]), .ZN(\Red_ToCheckInst_LFInst_35_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_35_LFInst_3_n2 ), .B(PermutationOutput[57]), 
        .ZN(Red_SignaltoCheck[143]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_3_U3  ( .A(PermutationOutput[58]), 
        .B(PermutationOutput[56]), .ZN(\Red_ToCheckInst_LFInst_35_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_36_LFInst_0_n2 ), .B(PermutationOutput[34]), 
        .ZN(Red_SignaltoCheck[144]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_0_U3  ( .A(PermutationOutput[35]), 
        .B(PermutationOutput[33]), .ZN(\Red_ToCheckInst_LFInst_36_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_36_LFInst_1_n2 ), .B(PermutationOutput[34]), 
        .ZN(Red_SignaltoCheck[145]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_1_U3  ( .A(PermutationOutput[35]), 
        .B(PermutationOutput[32]), .ZN(\Red_ToCheckInst_LFInst_36_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_36_LFInst_2_n2 ), .B(PermutationOutput[33]), 
        .ZN(Red_SignaltoCheck[146]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_2_U3  ( .A(PermutationOutput[35]), 
        .B(PermutationOutput[32]), .ZN(\Red_ToCheckInst_LFInst_36_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_36_LFInst_3_n2 ), .B(PermutationOutput[33]), 
        .ZN(Red_SignaltoCheck[147]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_3_U3  ( .A(PermutationOutput[34]), 
        .B(PermutationOutput[32]), .ZN(\Red_ToCheckInst_LFInst_36_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_37_LFInst_0_n2 ), .B(PermutationOutput[46]), 
        .ZN(Red_SignaltoCheck[148]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_0_U3  ( .A(PermutationOutput[47]), 
        .B(PermutationOutput[45]), .ZN(\Red_ToCheckInst_LFInst_37_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_37_LFInst_1_n2 ), .B(PermutationOutput[46]), 
        .ZN(Red_SignaltoCheck[149]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_1_U3  ( .A(PermutationOutput[47]), 
        .B(PermutationOutput[44]), .ZN(\Red_ToCheckInst_LFInst_37_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_37_LFInst_2_n2 ), .B(PermutationOutput[45]), 
        .ZN(Red_SignaltoCheck[150]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_2_U3  ( .A(PermutationOutput[47]), 
        .B(PermutationOutput[44]), .ZN(\Red_ToCheckInst_LFInst_37_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_37_LFInst_3_n2 ), .B(PermutationOutput[45]), 
        .ZN(Red_SignaltoCheck[151]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_3_U3  ( .A(PermutationOutput[46]), 
        .B(PermutationOutput[44]), .ZN(\Red_ToCheckInst_LFInst_37_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_38_LFInst_0_n2 ), .B(PermutationOutput[42]), 
        .ZN(Red_SignaltoCheck[152]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_0_U3  ( .A(PermutationOutput[43]), 
        .B(PermutationOutput[41]), .ZN(\Red_ToCheckInst_LFInst_38_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_38_LFInst_1_n2 ), .B(PermutationOutput[42]), 
        .ZN(Red_SignaltoCheck[153]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_1_U3  ( .A(PermutationOutput[43]), 
        .B(PermutationOutput[40]), .ZN(\Red_ToCheckInst_LFInst_38_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_38_LFInst_2_n2 ), .B(PermutationOutput[41]), 
        .ZN(Red_SignaltoCheck[154]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_2_U3  ( .A(PermutationOutput[43]), 
        .B(PermutationOutput[40]), .ZN(\Red_ToCheckInst_LFInst_38_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_38_LFInst_3_n2 ), .B(PermutationOutput[41]), 
        .ZN(Red_SignaltoCheck[155]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_3_U3  ( .A(PermutationOutput[42]), 
        .B(PermutationOutput[40]), .ZN(\Red_ToCheckInst_LFInst_38_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_39_LFInst_0_n2 ), .B(PermutationOutput[38]), 
        .ZN(Red_SignaltoCheck[156]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_0_U3  ( .A(PermutationOutput[39]), 
        .B(PermutationOutput[37]), .ZN(\Red_ToCheckInst_LFInst_39_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_39_LFInst_1_n2 ), .B(PermutationOutput[38]), 
        .ZN(Red_SignaltoCheck[157]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_1_U3  ( .A(PermutationOutput[39]), 
        .B(PermutationOutput[36]), .ZN(\Red_ToCheckInst_LFInst_39_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_39_LFInst_2_n2 ), .B(PermutationOutput[37]), 
        .ZN(Red_SignaltoCheck[158]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_2_U3  ( .A(PermutationOutput[39]), 
        .B(PermutationOutput[36]), .ZN(\Red_ToCheckInst_LFInst_39_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_39_LFInst_3_n2 ), .B(PermutationOutput[37]), 
        .ZN(Red_SignaltoCheck[159]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_3_U3  ( .A(PermutationOutput[38]), 
        .B(PermutationOutput[36]), .ZN(\Red_ToCheckInst_LFInst_39_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_40_LFInst_0_n2 ), .B(PermutationOutput[18]), 
        .ZN(Red_SignaltoCheck[160]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_0_U3  ( .A(PermutationOutput[19]), 
        .B(PermutationOutput[17]), .ZN(\Red_ToCheckInst_LFInst_40_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_40_LFInst_1_n2 ), .B(PermutationOutput[18]), 
        .ZN(Red_SignaltoCheck[161]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_1_U3  ( .A(PermutationOutput[19]), 
        .B(PermutationOutput[16]), .ZN(\Red_ToCheckInst_LFInst_40_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_40_LFInst_2_n2 ), .B(PermutationOutput[17]), 
        .ZN(Red_SignaltoCheck[162]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_2_U3  ( .A(PermutationOutput[19]), 
        .B(PermutationOutput[16]), .ZN(\Red_ToCheckInst_LFInst_40_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_40_LFInst_3_n2 ), .B(PermutationOutput[17]), 
        .ZN(Red_SignaltoCheck[163]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_3_U3  ( .A(PermutationOutput[18]), 
        .B(PermutationOutput[16]), .ZN(\Red_ToCheckInst_LFInst_40_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_41_LFInst_0_n2 ), .B(PermutationOutput[30]), 
        .ZN(Red_SignaltoCheck[164]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_0_U3  ( .A(PermutationOutput[31]), 
        .B(PermutationOutput[29]), .ZN(\Red_ToCheckInst_LFInst_41_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_41_LFInst_1_n2 ), .B(PermutationOutput[30]), 
        .ZN(Red_SignaltoCheck[165]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_1_U3  ( .A(PermutationOutput[31]), 
        .B(PermutationOutput[28]), .ZN(\Red_ToCheckInst_LFInst_41_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_41_LFInst_2_n2 ), .B(PermutationOutput[29]), 
        .ZN(Red_SignaltoCheck[166]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_2_U3  ( .A(PermutationOutput[31]), 
        .B(PermutationOutput[28]), .ZN(\Red_ToCheckInst_LFInst_41_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_41_LFInst_3_n2 ), .B(PermutationOutput[29]), 
        .ZN(Red_SignaltoCheck[167]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_3_U3  ( .A(PermutationOutput[30]), 
        .B(PermutationOutput[28]), .ZN(\Red_ToCheckInst_LFInst_41_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_42_LFInst_0_n2 ), .B(PermutationOutput[26]), 
        .ZN(Red_SignaltoCheck[168]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_0_U3  ( .A(PermutationOutput[27]), 
        .B(PermutationOutput[25]), .ZN(\Red_ToCheckInst_LFInst_42_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_42_LFInst_1_n2 ), .B(PermutationOutput[26]), 
        .ZN(Red_SignaltoCheck[169]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_1_U3  ( .A(PermutationOutput[27]), 
        .B(PermutationOutput[24]), .ZN(\Red_ToCheckInst_LFInst_42_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_42_LFInst_2_n2 ), .B(PermutationOutput[25]), 
        .ZN(Red_SignaltoCheck[170]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_2_U3  ( .A(PermutationOutput[27]), 
        .B(PermutationOutput[24]), .ZN(\Red_ToCheckInst_LFInst_42_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_42_LFInst_3_n2 ), .B(PermutationOutput[25]), 
        .ZN(Red_SignaltoCheck[171]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_3_U3  ( .A(PermutationOutput[26]), 
        .B(PermutationOutput[24]), .ZN(\Red_ToCheckInst_LFInst_42_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_43_LFInst_0_n2 ), .B(PermutationOutput[22]), 
        .ZN(Red_SignaltoCheck[172]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_0_U3  ( .A(PermutationOutput[23]), 
        .B(PermutationOutput[21]), .ZN(\Red_ToCheckInst_LFInst_43_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_43_LFInst_1_n2 ), .B(PermutationOutput[22]), 
        .ZN(Red_SignaltoCheck[173]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_1_U3  ( .A(PermutationOutput[23]), 
        .B(PermutationOutput[20]), .ZN(\Red_ToCheckInst_LFInst_43_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_43_LFInst_2_n2 ), .B(PermutationOutput[21]), 
        .ZN(Red_SignaltoCheck[174]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_2_U3  ( .A(PermutationOutput[23]), 
        .B(PermutationOutput[20]), .ZN(\Red_ToCheckInst_LFInst_43_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_43_LFInst_3_n2 ), .B(PermutationOutput[21]), 
        .ZN(Red_SignaltoCheck[175]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_3_U3  ( .A(PermutationOutput[22]), 
        .B(PermutationOutput[20]), .ZN(\Red_ToCheckInst_LFInst_43_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_44_LFInst_0_n2 ), .B(PermutationOutput[6]), 
        .ZN(Red_SignaltoCheck[176]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_0_U3  ( .A(PermutationOutput[7]), 
        .B(PermutationOutput[5]), .ZN(\Red_ToCheckInst_LFInst_44_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_44_LFInst_1_n2 ), .B(PermutationOutput[6]), 
        .ZN(Red_SignaltoCheck[177]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_1_U3  ( .A(PermutationOutput[7]), 
        .B(PermutationOutput[4]), .ZN(\Red_ToCheckInst_LFInst_44_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_44_LFInst_2_n2 ), .B(PermutationOutput[5]), 
        .ZN(Red_SignaltoCheck[178]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_2_U3  ( .A(PermutationOutput[7]), 
        .B(PermutationOutput[4]), .ZN(\Red_ToCheckInst_LFInst_44_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_44_LFInst_3_n2 ), .B(PermutationOutput[5]), 
        .ZN(Red_SignaltoCheck[179]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_3_U3  ( .A(PermutationOutput[6]), 
        .B(PermutationOutput[4]), .ZN(\Red_ToCheckInst_LFInst_44_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_45_LFInst_0_n2 ), .B(PermutationOutput[10]), 
        .ZN(Red_SignaltoCheck[180]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_0_U3  ( .A(PermutationOutput[11]), 
        .B(PermutationOutput[9]), .ZN(\Red_ToCheckInst_LFInst_45_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_45_LFInst_1_n2 ), .B(PermutationOutput[10]), 
        .ZN(Red_SignaltoCheck[181]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_1_U3  ( .A(PermutationOutput[11]), 
        .B(PermutationOutput[8]), .ZN(\Red_ToCheckInst_LFInst_45_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_45_LFInst_2_n2 ), .B(PermutationOutput[9]), 
        .ZN(Red_SignaltoCheck[182]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_2_U3  ( .A(PermutationOutput[11]), 
        .B(PermutationOutput[8]), .ZN(\Red_ToCheckInst_LFInst_45_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_45_LFInst_3_n2 ), .B(PermutationOutput[9]), 
        .ZN(Red_SignaltoCheck[183]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_3_U3  ( .A(PermutationOutput[10]), 
        .B(PermutationOutput[8]), .ZN(\Red_ToCheckInst_LFInst_45_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_46_LFInst_0_n2 ), .B(PermutationOutput[14]), 
        .ZN(Red_SignaltoCheck[184]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_0_U3  ( .A(PermutationOutput[15]), 
        .B(PermutationOutput[13]), .ZN(\Red_ToCheckInst_LFInst_46_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_46_LFInst_1_n2 ), .B(PermutationOutput[14]), 
        .ZN(Red_SignaltoCheck[185]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_1_U3  ( .A(PermutationOutput[15]), 
        .B(PermutationOutput[12]), .ZN(\Red_ToCheckInst_LFInst_46_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_46_LFInst_2_n2 ), .B(PermutationOutput[13]), 
        .ZN(Red_SignaltoCheck[186]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_2_U3  ( .A(PermutationOutput[15]), 
        .B(PermutationOutput[12]), .ZN(\Red_ToCheckInst_LFInst_46_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_46_LFInst_3_n2 ), .B(PermutationOutput[13]), 
        .ZN(Red_SignaltoCheck[187]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_3_U3  ( .A(PermutationOutput[14]), 
        .B(PermutationOutput[12]), .ZN(\Red_ToCheckInst_LFInst_46_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_47_LFInst_0_n2 ), .B(PermutationOutput[2]), 
        .ZN(Red_SignaltoCheck[188]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_0_U3  ( .A(PermutationOutput[3]), 
        .B(PermutationOutput[1]), .ZN(\Red_ToCheckInst_LFInst_47_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_47_LFInst_1_n2 ), .B(PermutationOutput[2]), 
        .ZN(Red_SignaltoCheck[189]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_1_U3  ( .A(PermutationOutput[3]), 
        .B(PermutationOutput[0]), .ZN(\Red_ToCheckInst_LFInst_47_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_47_LFInst_2_n2 ), .B(PermutationOutput[1]), 
        .ZN(Red_SignaltoCheck[190]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_2_U3  ( .A(PermutationOutput[3]), 
        .B(PermutationOutput[0]), .ZN(\Red_ToCheckInst_LFInst_47_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_47_LFInst_3_n2 ), .B(PermutationOutput[1]), 
        .ZN(Red_SignaltoCheck[191]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_3_U3  ( .A(PermutationOutput[2]), 
        .B(PermutationOutput[0]), .ZN(\Red_ToCheckInst_LFInst_47_LFInst_3_n2 )
         );
  NOR2_X1 \Check1_CheckInst_0_U95  ( .A1(\Check1_CheckInst_0_n94 ), .A2(
        \Check1_CheckInst_0_n93 ), .ZN(Error[0]) );
  NAND2_X1 \Check1_CheckInst_0_U94  ( .A1(\Check1_CheckInst_0_n92 ), .A2(
        \Check1_CheckInst_0_n91 ), .ZN(\Check1_CheckInst_0_n93 ) );
  NOR2_X1 \Check1_CheckInst_0_U93  ( .A1(\Check1_CheckInst_0_n90 ), .A2(
        \Check1_CheckInst_0_n89 ), .ZN(\Check1_CheckInst_0_n91 ) );
  NAND2_X1 \Check1_CheckInst_0_U92  ( .A1(\Check1_CheckInst_0_n88 ), .A2(
        \Check1_CheckInst_0_n87 ), .ZN(\Check1_CheckInst_0_n89 ) );
  NOR2_X1 \Check1_CheckInst_0_U91  ( .A1(\Check1_CheckInst_0_n86 ), .A2(
        \Check1_CheckInst_0_n85 ), .ZN(\Check1_CheckInst_0_n87 ) );
  NAND2_X1 \Check1_CheckInst_0_U90  ( .A1(\Check1_CheckInst_0_n84 ), .A2(
        \Check1_CheckInst_0_n83 ), .ZN(\Check1_CheckInst_0_n85 ) );
  NOR2_X1 \Check1_CheckInst_0_U89  ( .A1(\Check1_CheckInst_0_n82 ), .A2(
        \Check1_CheckInst_0_n81 ), .ZN(\Check1_CheckInst_0_n83 ) );
  NAND2_X1 \Check1_CheckInst_0_U88  ( .A1(\Check1_CheckInst_0_n80 ), .A2(
        \Check1_CheckInst_0_n79 ), .ZN(\Check1_CheckInst_0_n81 ) );
  XNOR2_X1 \Check1_CheckInst_0_U87  ( .A(Red_StateRegOutput[24]), .B(
        Red_SignaltoCheck[152]), .ZN(\Check1_CheckInst_0_n79 ) );
  XNOR2_X1 \Check1_CheckInst_0_U86  ( .A(Red_StateRegOutput[28]), .B(
        Red_SignaltoCheck[156]), .ZN(\Check1_CheckInst_0_n80 ) );
  NAND2_X1 \Check1_CheckInst_0_U85  ( .A1(\Check1_CheckInst_0_n78 ), .A2(
        \Check1_CheckInst_0_n77 ), .ZN(\Check1_CheckInst_0_n82 ) );
  XNOR2_X1 \Check1_CheckInst_0_U84  ( .A(Red_StateRegOutput[44]), .B(
        Red_SignaltoCheck[172]), .ZN(\Check1_CheckInst_0_n77 ) );
  XNOR2_X1 \Check1_CheckInst_0_U83  ( .A(Red_StateRegOutput[36]), .B(
        Red_SignaltoCheck[164]), .ZN(\Check1_CheckInst_0_n78 ) );
  NOR2_X1 \Check1_CheckInst_0_U82  ( .A1(\Check1_CheckInst_0_n76 ), .A2(
        \Check1_CheckInst_0_n75 ), .ZN(\Check1_CheckInst_0_n84 ) );
  NAND2_X1 \Check1_CheckInst_0_U81  ( .A1(\Check1_CheckInst_0_n74 ), .A2(
        \Check1_CheckInst_0_n73 ), .ZN(\Check1_CheckInst_0_n75 ) );
  XNOR2_X1 \Check1_CheckInst_0_U80  ( .A(Red_StateRegOutput[20]), .B(
        Red_SignaltoCheck[148]), .ZN(\Check1_CheckInst_0_n73 ) );
  XNOR2_X1 \Check1_CheckInst_0_U79  ( .A(Red_StateRegOutput[12]), .B(
        Red_SignaltoCheck[140]), .ZN(\Check1_CheckInst_0_n74 ) );
  NAND2_X1 \Check1_CheckInst_0_U78  ( .A1(\Check1_CheckInst_0_n72 ), .A2(
        \Check1_CheckInst_0_n71 ), .ZN(\Check1_CheckInst_0_n76 ) );
  XNOR2_X1 \Check1_CheckInst_0_U77  ( .A(Red_StateRegOutput[16]), .B(
        Red_SignaltoCheck[144]), .ZN(\Check1_CheckInst_0_n71 ) );
  XNOR2_X1 \Check1_CheckInst_0_U76  ( .A(Red_StateRegOutput[32]), .B(
        Red_SignaltoCheck[160]), .ZN(\Check1_CheckInst_0_n72 ) );
  NAND2_X1 \Check1_CheckInst_0_U75  ( .A1(\Check1_CheckInst_0_n70 ), .A2(
        \Check1_CheckInst_0_n69 ), .ZN(\Check1_CheckInst_0_n86 ) );
  NOR2_X1 \Check1_CheckInst_0_U74  ( .A1(\Check1_CheckInst_0_n68 ), .A2(
        \Check1_CheckInst_0_n67 ), .ZN(\Check1_CheckInst_0_n69 ) );
  XOR2_X1 \Check1_CheckInst_0_U73  ( .A(Red_AddRoundKeyOutput[24]), .B(
        Red_SignaltoCheck[24]), .Z(\Check1_CheckInst_0_n67 ) );
  XOR2_X1 \Check1_CheckInst_0_U72  ( .A(Red_AddRoundKeyOutput[40]), .B(
        Red_SignaltoCheck[40]), .Z(\Check1_CheckInst_0_n68 ) );
  NOR2_X1 \Check1_CheckInst_0_U71  ( .A1(\Check1_CheckInst_0_n66 ), .A2(
        \Check1_CheckInst_0_n65 ), .ZN(\Check1_CheckInst_0_n70 ) );
  XOR2_X1 \Check1_CheckInst_0_U70  ( .A(Red_AddRoundKeyOutput[32]), .B(
        Red_SignaltoCheck[32]), .Z(\Check1_CheckInst_0_n65 ) );
  XOR2_X1 \Check1_CheckInst_0_U69  ( .A(Red_AddRoundKeyOutput[36]), .B(
        Red_SignaltoCheck[36]), .Z(\Check1_CheckInst_0_n66 ) );
  NOR2_X1 \Check1_CheckInst_0_U68  ( .A1(\Check1_CheckInst_0_n64 ), .A2(
        \Check1_CheckInst_0_n63 ), .ZN(\Check1_CheckInst_0_n88 ) );
  NAND2_X1 \Check1_CheckInst_0_U67  ( .A1(\Check1_CheckInst_0_n62 ), .A2(
        \Check1_CheckInst_0_n61 ), .ZN(\Check1_CheckInst_0_n63 ) );
  XNOR2_X1 \Check1_CheckInst_0_U66  ( .A(Red_AddRoundKeyOutput[8]), .B(
        Red_SignaltoCheck[8]), .ZN(\Check1_CheckInst_0_n61 ) );
  XNOR2_X1 \Check1_CheckInst_0_U65  ( .A(Red_AddRoundKeyOutput[12]), .B(
        Red_SignaltoCheck[12]), .ZN(\Check1_CheckInst_0_n62 ) );
  NAND2_X1 \Check1_CheckInst_0_U64  ( .A1(\Check1_CheckInst_0_n60 ), .A2(
        \Check1_CheckInst_0_n59 ), .ZN(\Check1_CheckInst_0_n64 ) );
  XNOR2_X1 \Check1_CheckInst_0_U63  ( .A(Red_AddRoundKeyOutput[28]), .B(
        Red_SignaltoCheck[28]), .ZN(\Check1_CheckInst_0_n59 ) );
  XNOR2_X1 \Check1_CheckInst_0_U62  ( .A(Red_AddRoundKeyOutput[20]), .B(
        Red_SignaltoCheck[20]), .ZN(\Check1_CheckInst_0_n60 ) );
  NAND2_X1 \Check1_CheckInst_0_U61  ( .A1(\Check1_CheckInst_0_n58 ), .A2(
        \Check1_CheckInst_0_n57 ), .ZN(\Check1_CheckInst_0_n90 ) );
  NOR2_X1 \Check1_CheckInst_0_U60  ( .A1(\Check1_CheckInst_0_n56 ), .A2(
        \Check1_CheckInst_0_n55 ), .ZN(\Check1_CheckInst_0_n57 ) );
  NAND2_X1 \Check1_CheckInst_0_U59  ( .A1(\Check1_CheckInst_0_n54 ), .A2(
        \Check1_CheckInst_0_n53 ), .ZN(\Check1_CheckInst_0_n55 ) );
  NOR2_X1 \Check1_CheckInst_0_U58  ( .A1(\Check1_CheckInst_0_n52 ), .A2(
        \Check1_CheckInst_0_n51 ), .ZN(\Check1_CheckInst_0_n53 ) );
  NAND2_X1 \Check1_CheckInst_0_U57  ( .A1(\Check1_CheckInst_0_n50 ), .A2(
        \Check1_CheckInst_0_n49 ), .ZN(\Check1_CheckInst_0_n51 ) );
  XNOR2_X1 \Check1_CheckInst_0_U56  ( .A(Red_StateRegOutput[60]), .B(
        Red_SignaltoCheck[188]), .ZN(\Check1_CheckInst_0_n49 ) );
  XNOR2_X1 \Check1_CheckInst_0_U55  ( .A(Red_SignaltoCheck[4]), .B(
        Red_AddRoundKeyOutput[4]), .ZN(\Check1_CheckInst_0_n50 ) );
  NAND2_X1 \Check1_CheckInst_0_U54  ( .A1(\Check1_CheckInst_0_n48 ), .A2(
        \Check1_CheckInst_0_n47 ), .ZN(\Check1_CheckInst_0_n52 ) );
  XNOR2_X1 \Check1_CheckInst_0_U53  ( .A(Red_AddRoundKeyOutput[0]), .B(
        Red_SignaltoCheck[0]), .ZN(\Check1_CheckInst_0_n47 ) );
  XNOR2_X1 \Check1_CheckInst_0_U52  ( .A(Red_AddRoundKeyOutput[16]), .B(
        Red_SignaltoCheck[16]), .ZN(\Check1_CheckInst_0_n48 ) );
  NOR2_X1 \Check1_CheckInst_0_U51  ( .A1(\Check1_CheckInst_0_n46 ), .A2(
        \Check1_CheckInst_0_n45 ), .ZN(\Check1_CheckInst_0_n54 ) );
  NAND2_X1 \Check1_CheckInst_0_U50  ( .A1(\Check1_CheckInst_0_n44 ), .A2(
        \Check1_CheckInst_0_n43 ), .ZN(\Check1_CheckInst_0_n45 ) );
  XNOR2_X1 \Check1_CheckInst_0_U49  ( .A(Red_Feedback[8]), .B(
        Red_SignaltoCheck[72]), .ZN(\Check1_CheckInst_0_n43 ) );
  XNOR2_X1 \Check1_CheckInst_0_U48  ( .A(Red_Feedback[24]), .B(
        Red_SignaltoCheck[88]), .ZN(\Check1_CheckInst_0_n44 ) );
  NAND2_X1 \Check1_CheckInst_0_U47  ( .A1(\Check1_CheckInst_0_n42 ), .A2(
        \Check1_CheckInst_0_n41 ), .ZN(\Check1_CheckInst_0_n46 ) );
  XNOR2_X1 \Check1_CheckInst_0_U46  ( .A(Red_Feedback[16]), .B(
        Red_SignaltoCheck[80]), .ZN(\Check1_CheckInst_0_n41 ) );
  XNOR2_X1 \Check1_CheckInst_0_U45  ( .A(Red_Feedback[20]), .B(
        Red_SignaltoCheck[84]), .ZN(\Check1_CheckInst_0_n42 ) );
  NAND2_X1 \Check1_CheckInst_0_U44  ( .A1(\Check1_CheckInst_0_n40 ), .A2(
        \Check1_CheckInst_0_n39 ), .ZN(\Check1_CheckInst_0_n56 ) );
  NOR2_X1 \Check1_CheckInst_0_U43  ( .A1(\Check1_CheckInst_0_n38 ), .A2(
        \Check1_CheckInst_0_n37 ), .ZN(\Check1_CheckInst_0_n39 ) );
  XOR2_X1 \Check1_CheckInst_0_U42  ( .A(Red_AddRoundKeyOutput[56]), .B(
        Red_SignaltoCheck[56]), .Z(\Check1_CheckInst_0_n37 ) );
  XOR2_X1 \Check1_CheckInst_0_U41  ( .A(Red_AddRoundKeyOutput[60]), .B(
        Red_SignaltoCheck[60]), .Z(\Check1_CheckInst_0_n38 ) );
  NOR2_X1 \Check1_CheckInst_0_U40  ( .A1(\Check1_CheckInst_0_n36 ), .A2(
        \Check1_CheckInst_0_n35 ), .ZN(\Check1_CheckInst_0_n40 ) );
  XOR2_X1 \Check1_CheckInst_0_U39  ( .A(Red_Feedback[12]), .B(
        Red_SignaltoCheck[76]), .Z(\Check1_CheckInst_0_n35 ) );
  XOR2_X1 \Check1_CheckInst_0_U38  ( .A(Red_Feedback[4]), .B(
        Red_SignaltoCheck[68]), .Z(\Check1_CheckInst_0_n36 ) );
  NOR2_X1 \Check1_CheckInst_0_U37  ( .A1(\Check1_CheckInst_0_n34 ), .A2(
        \Check1_CheckInst_0_n33 ), .ZN(\Check1_CheckInst_0_n58 ) );
  NAND2_X1 \Check1_CheckInst_0_U36  ( .A1(\Check1_CheckInst_0_n32 ), .A2(
        \Check1_CheckInst_0_n31 ), .ZN(\Check1_CheckInst_0_n33 ) );
  XNOR2_X1 \Check1_CheckInst_0_U35  ( .A(Red_AddRoundKeyOutput[52]), .B(
        Red_SignaltoCheck[52]), .ZN(\Check1_CheckInst_0_n31 ) );
  XNOR2_X1 \Check1_CheckInst_0_U34  ( .A(Red_AddRoundKeyOutput[44]), .B(
        Red_SignaltoCheck[44]), .ZN(\Check1_CheckInst_0_n32 ) );
  NAND2_X1 \Check1_CheckInst_0_U33  ( .A1(\Check1_CheckInst_0_n30 ), .A2(
        \Check1_CheckInst_0_n29 ), .ZN(\Check1_CheckInst_0_n34 ) );
  XNOR2_X1 \Check1_CheckInst_0_U32  ( .A(Red_AddRoundKeyOutput[48]), .B(
        Red_SignaltoCheck[48]), .ZN(\Check1_CheckInst_0_n29 ) );
  XNOR2_X1 \Check1_CheckInst_0_U31  ( .A(Red_Feedback[0]), .B(
        Red_SignaltoCheck[64]), .ZN(\Check1_CheckInst_0_n30 ) );
  NOR2_X1 \Check1_CheckInst_0_U30  ( .A1(\Check1_CheckInst_0_n28 ), .A2(
        \Check1_CheckInst_0_n27 ), .ZN(\Check1_CheckInst_0_n92 ) );
  NAND2_X1 \Check1_CheckInst_0_U29  ( .A1(\Check1_CheckInst_0_n26 ), .A2(
        \Check1_CheckInst_0_n25 ), .ZN(\Check1_CheckInst_0_n27 ) );
  NOR2_X1 \Check1_CheckInst_0_U28  ( .A1(\Check1_CheckInst_0_n24 ), .A2(
        \Check1_CheckInst_0_n23 ), .ZN(\Check1_CheckInst_0_n25 ) );
  NAND2_X1 \Check1_CheckInst_0_U27  ( .A1(\Check1_CheckInst_0_n22 ), .A2(
        \Check1_CheckInst_0_n21 ), .ZN(\Check1_CheckInst_0_n23 ) );
  XNOR2_X1 \Check1_CheckInst_0_U26  ( .A(Red_StateRegOutput[0]), .B(
        Red_SignaltoCheck[128]), .ZN(\Check1_CheckInst_0_n21 ) );
  XNOR2_X1 \Check1_CheckInst_0_U25  ( .A(Red_StateRegOutput[4]), .B(
        Red_SignaltoCheck[132]), .ZN(\Check1_CheckInst_0_n22 ) );
  NAND2_X1 \Check1_CheckInst_0_U24  ( .A1(\Check1_CheckInst_0_n20 ), .A2(
        \Check1_CheckInst_0_n19 ), .ZN(\Check1_CheckInst_0_n24 ) );
  XNOR2_X1 \Check1_CheckInst_0_U23  ( .A(Red_Feedback[56]), .B(
        Red_SignaltoCheck[120]), .ZN(\Check1_CheckInst_0_n19 ) );
  XNOR2_X1 \Check1_CheckInst_0_U22  ( .A(Red_StateRegOutput[8]), .B(
        Red_SignaltoCheck[136]), .ZN(\Check1_CheckInst_0_n20 ) );
  NOR2_X1 \Check1_CheckInst_0_U21  ( .A1(\Check1_CheckInst_0_n18 ), .A2(
        \Check1_CheckInst_0_n17 ), .ZN(\Check1_CheckInst_0_n26 ) );
  XOR2_X1 \Check1_CheckInst_0_U20  ( .A(Red_Feedback[60]), .B(
        Red_SignaltoCheck[124]), .Z(\Check1_CheckInst_0_n17 ) );
  XOR2_X1 \Check1_CheckInst_0_U19  ( .A(Red_Feedback[52]), .B(
        Red_SignaltoCheck[116]), .Z(\Check1_CheckInst_0_n18 ) );
  NAND2_X1 \Check1_CheckInst_0_U18  ( .A1(\Check1_CheckInst_0_n16 ), .A2(
        \Check1_CheckInst_0_n15 ), .ZN(\Check1_CheckInst_0_n28 ) );
  XNOR2_X1 \Check1_CheckInst_0_U17  ( .A(Red_Feedback[40]), .B(
        Red_SignaltoCheck[104]), .ZN(\Check1_CheckInst_0_n15 ) );
  XNOR2_X1 \Check1_CheckInst_0_U16  ( .A(Red_Feedback[44]), .B(
        Red_SignaltoCheck[108]), .ZN(\Check1_CheckInst_0_n16 ) );
  NAND2_X1 \Check1_CheckInst_0_U15  ( .A1(\Check1_CheckInst_0_n14 ), .A2(
        \Check1_CheckInst_0_n13 ), .ZN(\Check1_CheckInst_0_n94 ) );
  NOR2_X1 \Check1_CheckInst_0_U14  ( .A1(\Check1_CheckInst_0_n12 ), .A2(
        \Check1_CheckInst_0_n11 ), .ZN(\Check1_CheckInst_0_n13 ) );
  NAND2_X1 \Check1_CheckInst_0_U13  ( .A1(\Check1_CheckInst_0_n10 ), .A2(
        \Check1_CheckInst_0_n9 ), .ZN(\Check1_CheckInst_0_n11 ) );
  NOR2_X1 \Check1_CheckInst_0_U12  ( .A1(\Check1_CheckInst_0_n8 ), .A2(
        \Check1_CheckInst_0_n7 ), .ZN(\Check1_CheckInst_0_n9 ) );
  XOR2_X1 \Check1_CheckInst_0_U11  ( .A(Red_Feedback[32]), .B(
        Red_SignaltoCheck[96]), .Z(\Check1_CheckInst_0_n7 ) );
  XOR2_X1 \Check1_CheckInst_0_U10  ( .A(Red_Feedback[48]), .B(
        Red_SignaltoCheck[112]), .Z(\Check1_CheckInst_0_n8 ) );
  NOR2_X1 \Check1_CheckInst_0_U9  ( .A1(\Check1_CheckInst_0_n6 ), .A2(
        \Check1_CheckInst_0_n5 ), .ZN(\Check1_CheckInst_0_n10 ) );
  XOR2_X1 \Check1_CheckInst_0_U8  ( .A(Red_Feedback[36]), .B(
        Red_SignaltoCheck[100]), .Z(\Check1_CheckInst_0_n5 ) );
  XOR2_X1 \Check1_CheckInst_0_U7  ( .A(Red_Feedback[28]), .B(
        Red_SignaltoCheck[92]), .Z(\Check1_CheckInst_0_n6 ) );
  NAND2_X1 \Check1_CheckInst_0_U6  ( .A1(\Check1_CheckInst_0_n4 ), .A2(
        \Check1_CheckInst_0_n3 ), .ZN(\Check1_CheckInst_0_n12 ) );
  XNOR2_X1 \Check1_CheckInst_0_U5  ( .A(Red_StateRegOutput[48]), .B(
        Red_SignaltoCheck[176]), .ZN(\Check1_CheckInst_0_n3 ) );
  XNOR2_X1 \Check1_CheckInst_0_U4  ( .A(Red_StateRegOutput[52]), .B(
        Red_SignaltoCheck[180]), .ZN(\Check1_CheckInst_0_n4 ) );
  NOR2_X1 \Check1_CheckInst_0_U3  ( .A1(\Check1_CheckInst_0_n2 ), .A2(
        \Check1_CheckInst_0_n1 ), .ZN(\Check1_CheckInst_0_n14 ) );
  XOR2_X1 \Check1_CheckInst_0_U2  ( .A(Red_StateRegOutput[40]), .B(
        Red_SignaltoCheck[168]), .Z(\Check1_CheckInst_0_n1 ) );
  XOR2_X1 \Check1_CheckInst_0_U1  ( .A(Red_StateRegOutput[56]), .B(
        Red_SignaltoCheck[184]), .Z(\Check1_CheckInst_0_n2 ) );
  NOR2_X1 \Check1_CheckInst_1_U95  ( .A1(\Check1_CheckInst_1_n96 ), .A2(
        \Check1_CheckInst_1_n95 ), .ZN(Error[1]) );
  NAND2_X1 \Check1_CheckInst_1_U94  ( .A1(\Check1_CheckInst_1_n94 ), .A2(
        \Check1_CheckInst_1_n93 ), .ZN(\Check1_CheckInst_1_n95 ) );
  NOR2_X1 \Check1_CheckInst_1_U93  ( .A1(\Check1_CheckInst_1_n92 ), .A2(
        \Check1_CheckInst_1_n91 ), .ZN(\Check1_CheckInst_1_n93 ) );
  NAND2_X1 \Check1_CheckInst_1_U92  ( .A1(\Check1_CheckInst_1_n90 ), .A2(
        \Check1_CheckInst_1_n89 ), .ZN(\Check1_CheckInst_1_n91 ) );
  NOR2_X1 \Check1_CheckInst_1_U91  ( .A1(\Check1_CheckInst_1_n88 ), .A2(
        \Check1_CheckInst_1_n87 ), .ZN(\Check1_CheckInst_1_n89 ) );
  NAND2_X1 \Check1_CheckInst_1_U90  ( .A1(\Check1_CheckInst_1_n86 ), .A2(
        \Check1_CheckInst_1_n85 ), .ZN(\Check1_CheckInst_1_n87 ) );
  NOR2_X1 \Check1_CheckInst_1_U89  ( .A1(\Check1_CheckInst_1_n84 ), .A2(
        \Check1_CheckInst_1_n83 ), .ZN(\Check1_CheckInst_1_n85 ) );
  NAND2_X1 \Check1_CheckInst_1_U88  ( .A1(\Check1_CheckInst_1_n82 ), .A2(
        \Check1_CheckInst_1_n81 ), .ZN(\Check1_CheckInst_1_n83 ) );
  XNOR2_X1 \Check1_CheckInst_1_U87  ( .A(Red_StateRegOutput[25]), .B(
        Red_SignaltoCheck[153]), .ZN(\Check1_CheckInst_1_n81 ) );
  XNOR2_X1 \Check1_CheckInst_1_U86  ( .A(Red_StateRegOutput[29]), .B(
        Red_SignaltoCheck[157]), .ZN(\Check1_CheckInst_1_n82 ) );
  NAND2_X1 \Check1_CheckInst_1_U85  ( .A1(\Check1_CheckInst_1_n80 ), .A2(
        \Check1_CheckInst_1_n79 ), .ZN(\Check1_CheckInst_1_n84 ) );
  XNOR2_X1 \Check1_CheckInst_1_U84  ( .A(Red_StateRegOutput[45]), .B(
        Red_SignaltoCheck[173]), .ZN(\Check1_CheckInst_1_n79 ) );
  XNOR2_X1 \Check1_CheckInst_1_U83  ( .A(Red_StateRegOutput[37]), .B(
        Red_SignaltoCheck[165]), .ZN(\Check1_CheckInst_1_n80 ) );
  NOR2_X1 \Check1_CheckInst_1_U82  ( .A1(\Check1_CheckInst_1_n78 ), .A2(
        \Check1_CheckInst_1_n77 ), .ZN(\Check1_CheckInst_1_n86 ) );
  NAND2_X1 \Check1_CheckInst_1_U81  ( .A1(\Check1_CheckInst_1_n76 ), .A2(
        \Check1_CheckInst_1_n75 ), .ZN(\Check1_CheckInst_1_n77 ) );
  XNOR2_X1 \Check1_CheckInst_1_U80  ( .A(Red_StateRegOutput[21]), .B(
        Red_SignaltoCheck[149]), .ZN(\Check1_CheckInst_1_n75 ) );
  XNOR2_X1 \Check1_CheckInst_1_U79  ( .A(Red_StateRegOutput[13]), .B(
        Red_SignaltoCheck[141]), .ZN(\Check1_CheckInst_1_n76 ) );
  NAND2_X1 \Check1_CheckInst_1_U78  ( .A1(\Check1_CheckInst_1_n74 ), .A2(
        \Check1_CheckInst_1_n73 ), .ZN(\Check1_CheckInst_1_n78 ) );
  XNOR2_X1 \Check1_CheckInst_1_U77  ( .A(Red_StateRegOutput[17]), .B(
        Red_SignaltoCheck[145]), .ZN(\Check1_CheckInst_1_n73 ) );
  XNOR2_X1 \Check1_CheckInst_1_U76  ( .A(Red_StateRegOutput[33]), .B(
        Red_SignaltoCheck[161]), .ZN(\Check1_CheckInst_1_n74 ) );
  NAND2_X1 \Check1_CheckInst_1_U75  ( .A1(\Check1_CheckInst_1_n72 ), .A2(
        \Check1_CheckInst_1_n71 ), .ZN(\Check1_CheckInst_1_n88 ) );
  NOR2_X1 \Check1_CheckInst_1_U74  ( .A1(\Check1_CheckInst_1_n70 ), .A2(
        \Check1_CheckInst_1_n69 ), .ZN(\Check1_CheckInst_1_n71 ) );
  XOR2_X1 \Check1_CheckInst_1_U73  ( .A(Red_AddRoundKeyOutput[25]), .B(
        Red_SignaltoCheck[25]), .Z(\Check1_CheckInst_1_n69 ) );
  XOR2_X1 \Check1_CheckInst_1_U72  ( .A(Red_AddRoundKeyOutput[41]), .B(
        Red_SignaltoCheck[41]), .Z(\Check1_CheckInst_1_n70 ) );
  NOR2_X1 \Check1_CheckInst_1_U71  ( .A1(\Check1_CheckInst_1_n68 ), .A2(
        \Check1_CheckInst_1_n67 ), .ZN(\Check1_CheckInst_1_n72 ) );
  XOR2_X1 \Check1_CheckInst_1_U70  ( .A(Red_AddRoundKeyOutput[33]), .B(
        Red_SignaltoCheck[33]), .Z(\Check1_CheckInst_1_n67 ) );
  XOR2_X1 \Check1_CheckInst_1_U69  ( .A(Red_AddRoundKeyOutput[37]), .B(
        Red_SignaltoCheck[37]), .Z(\Check1_CheckInst_1_n68 ) );
  NOR2_X1 \Check1_CheckInst_1_U68  ( .A1(\Check1_CheckInst_1_n66 ), .A2(
        \Check1_CheckInst_1_n65 ), .ZN(\Check1_CheckInst_1_n90 ) );
  NAND2_X1 \Check1_CheckInst_1_U67  ( .A1(\Check1_CheckInst_1_n64 ), .A2(
        \Check1_CheckInst_1_n63 ), .ZN(\Check1_CheckInst_1_n65 ) );
  XNOR2_X1 \Check1_CheckInst_1_U66  ( .A(Red_AddRoundKeyOutput[9]), .B(
        Red_SignaltoCheck[9]), .ZN(\Check1_CheckInst_1_n63 ) );
  XNOR2_X1 \Check1_CheckInst_1_U65  ( .A(Red_AddRoundKeyOutput[13]), .B(
        Red_SignaltoCheck[13]), .ZN(\Check1_CheckInst_1_n64 ) );
  NAND2_X1 \Check1_CheckInst_1_U64  ( .A1(\Check1_CheckInst_1_n62 ), .A2(
        \Check1_CheckInst_1_n61 ), .ZN(\Check1_CheckInst_1_n66 ) );
  XNOR2_X1 \Check1_CheckInst_1_U63  ( .A(Red_AddRoundKeyOutput[29]), .B(
        Red_SignaltoCheck[29]), .ZN(\Check1_CheckInst_1_n61 ) );
  XNOR2_X1 \Check1_CheckInst_1_U62  ( .A(Red_AddRoundKeyOutput[21]), .B(
        Red_SignaltoCheck[21]), .ZN(\Check1_CheckInst_1_n62 ) );
  NAND2_X1 \Check1_CheckInst_1_U61  ( .A1(\Check1_CheckInst_1_n60 ), .A2(
        \Check1_CheckInst_1_n59 ), .ZN(\Check1_CheckInst_1_n92 ) );
  NOR2_X1 \Check1_CheckInst_1_U60  ( .A1(\Check1_CheckInst_1_n58 ), .A2(
        \Check1_CheckInst_1_n57 ), .ZN(\Check1_CheckInst_1_n59 ) );
  NAND2_X1 \Check1_CheckInst_1_U59  ( .A1(\Check1_CheckInst_1_n56 ), .A2(
        \Check1_CheckInst_1_n55 ), .ZN(\Check1_CheckInst_1_n57 ) );
  NOR2_X1 \Check1_CheckInst_1_U58  ( .A1(\Check1_CheckInst_1_n54 ), .A2(
        \Check1_CheckInst_1_n53 ), .ZN(\Check1_CheckInst_1_n55 ) );
  NAND2_X1 \Check1_CheckInst_1_U57  ( .A1(\Check1_CheckInst_1_n52 ), .A2(
        \Check1_CheckInst_1_n51 ), .ZN(\Check1_CheckInst_1_n53 ) );
  XNOR2_X1 \Check1_CheckInst_1_U56  ( .A(Red_StateRegOutput[61]), .B(
        Red_SignaltoCheck[189]), .ZN(\Check1_CheckInst_1_n51 ) );
  XNOR2_X1 \Check1_CheckInst_1_U55  ( .A(Red_SignaltoCheck[5]), .B(
        Red_AddRoundKeyOutput[5]), .ZN(\Check1_CheckInst_1_n52 ) );
  NAND2_X1 \Check1_CheckInst_1_U54  ( .A1(\Check1_CheckInst_1_n50 ), .A2(
        \Check1_CheckInst_1_n49 ), .ZN(\Check1_CheckInst_1_n54 ) );
  XNOR2_X1 \Check1_CheckInst_1_U53  ( .A(Red_AddRoundKeyOutput[1]), .B(
        Red_SignaltoCheck[1]), .ZN(\Check1_CheckInst_1_n49 ) );
  XNOR2_X1 \Check1_CheckInst_1_U52  ( .A(Red_AddRoundKeyOutput[17]), .B(
        Red_SignaltoCheck[17]), .ZN(\Check1_CheckInst_1_n50 ) );
  NOR2_X1 \Check1_CheckInst_1_U51  ( .A1(\Check1_CheckInst_1_n48 ), .A2(
        \Check1_CheckInst_1_n47 ), .ZN(\Check1_CheckInst_1_n56 ) );
  NAND2_X1 \Check1_CheckInst_1_U50  ( .A1(\Check1_CheckInst_1_n46 ), .A2(
        \Check1_CheckInst_1_n45 ), .ZN(\Check1_CheckInst_1_n47 ) );
  XNOR2_X1 \Check1_CheckInst_1_U49  ( .A(Red_Feedback[9]), .B(
        Red_SignaltoCheck[73]), .ZN(\Check1_CheckInst_1_n45 ) );
  XNOR2_X1 \Check1_CheckInst_1_U48  ( .A(Red_Feedback[25]), .B(
        Red_SignaltoCheck[89]), .ZN(\Check1_CheckInst_1_n46 ) );
  NAND2_X1 \Check1_CheckInst_1_U47  ( .A1(\Check1_CheckInst_1_n44 ), .A2(
        \Check1_CheckInst_1_n43 ), .ZN(\Check1_CheckInst_1_n48 ) );
  XNOR2_X1 \Check1_CheckInst_1_U46  ( .A(Red_Feedback[17]), .B(
        Red_SignaltoCheck[81]), .ZN(\Check1_CheckInst_1_n43 ) );
  XNOR2_X1 \Check1_CheckInst_1_U45  ( .A(Red_Feedback[21]), .B(
        Red_SignaltoCheck[85]), .ZN(\Check1_CheckInst_1_n44 ) );
  NAND2_X1 \Check1_CheckInst_1_U44  ( .A1(\Check1_CheckInst_1_n42 ), .A2(
        \Check1_CheckInst_1_n41 ), .ZN(\Check1_CheckInst_1_n58 ) );
  NOR2_X1 \Check1_CheckInst_1_U43  ( .A1(\Check1_CheckInst_1_n40 ), .A2(
        \Check1_CheckInst_1_n39 ), .ZN(\Check1_CheckInst_1_n41 ) );
  XOR2_X1 \Check1_CheckInst_1_U42  ( .A(Red_AddRoundKeyOutput[57]), .B(
        Red_SignaltoCheck[57]), .Z(\Check1_CheckInst_1_n39 ) );
  XOR2_X1 \Check1_CheckInst_1_U41  ( .A(Red_AddRoundKeyOutput[61]), .B(
        Red_SignaltoCheck[61]), .Z(\Check1_CheckInst_1_n40 ) );
  NOR2_X1 \Check1_CheckInst_1_U40  ( .A1(\Check1_CheckInst_1_n38 ), .A2(
        \Check1_CheckInst_1_n37 ), .ZN(\Check1_CheckInst_1_n42 ) );
  XOR2_X1 \Check1_CheckInst_1_U39  ( .A(Red_Feedback[13]), .B(
        Red_SignaltoCheck[77]), .Z(\Check1_CheckInst_1_n37 ) );
  XOR2_X1 \Check1_CheckInst_1_U38  ( .A(Red_Feedback[5]), .B(
        Red_SignaltoCheck[69]), .Z(\Check1_CheckInst_1_n38 ) );
  NOR2_X1 \Check1_CheckInst_1_U37  ( .A1(\Check1_CheckInst_1_n36 ), .A2(
        \Check1_CheckInst_1_n35 ), .ZN(\Check1_CheckInst_1_n60 ) );
  NAND2_X1 \Check1_CheckInst_1_U36  ( .A1(\Check1_CheckInst_1_n34 ), .A2(
        \Check1_CheckInst_1_n33 ), .ZN(\Check1_CheckInst_1_n35 ) );
  XNOR2_X1 \Check1_CheckInst_1_U35  ( .A(Red_AddRoundKeyOutput[53]), .B(
        Red_SignaltoCheck[53]), .ZN(\Check1_CheckInst_1_n33 ) );
  XNOR2_X1 \Check1_CheckInst_1_U34  ( .A(Red_AddRoundKeyOutput[45]), .B(
        Red_SignaltoCheck[45]), .ZN(\Check1_CheckInst_1_n34 ) );
  NAND2_X1 \Check1_CheckInst_1_U33  ( .A1(\Check1_CheckInst_1_n32 ), .A2(
        \Check1_CheckInst_1_n31 ), .ZN(\Check1_CheckInst_1_n36 ) );
  XNOR2_X1 \Check1_CheckInst_1_U32  ( .A(Red_AddRoundKeyOutput[49]), .B(
        Red_SignaltoCheck[49]), .ZN(\Check1_CheckInst_1_n31 ) );
  XNOR2_X1 \Check1_CheckInst_1_U31  ( .A(Red_Feedback[1]), .B(
        Red_SignaltoCheck[65]), .ZN(\Check1_CheckInst_1_n32 ) );
  NOR2_X1 \Check1_CheckInst_1_U30  ( .A1(\Check1_CheckInst_1_n30 ), .A2(
        \Check1_CheckInst_1_n29 ), .ZN(\Check1_CheckInst_1_n94 ) );
  NAND2_X1 \Check1_CheckInst_1_U29  ( .A1(\Check1_CheckInst_1_n28 ), .A2(
        \Check1_CheckInst_1_n27 ), .ZN(\Check1_CheckInst_1_n29 ) );
  NOR2_X1 \Check1_CheckInst_1_U28  ( .A1(\Check1_CheckInst_1_n26 ), .A2(
        \Check1_CheckInst_1_n25 ), .ZN(\Check1_CheckInst_1_n27 ) );
  NAND2_X1 \Check1_CheckInst_1_U27  ( .A1(\Check1_CheckInst_1_n24 ), .A2(
        \Check1_CheckInst_1_n23 ), .ZN(\Check1_CheckInst_1_n25 ) );
  XNOR2_X1 \Check1_CheckInst_1_U26  ( .A(Red_StateRegOutput[1]), .B(
        Red_SignaltoCheck[129]), .ZN(\Check1_CheckInst_1_n23 ) );
  XNOR2_X1 \Check1_CheckInst_1_U25  ( .A(Red_StateRegOutput[5]), .B(
        Red_SignaltoCheck[133]), .ZN(\Check1_CheckInst_1_n24 ) );
  NAND2_X1 \Check1_CheckInst_1_U24  ( .A1(\Check1_CheckInst_1_n22 ), .A2(
        \Check1_CheckInst_1_n21 ), .ZN(\Check1_CheckInst_1_n26 ) );
  XNOR2_X1 \Check1_CheckInst_1_U23  ( .A(Red_Feedback[57]), .B(
        Red_SignaltoCheck[121]), .ZN(\Check1_CheckInst_1_n21 ) );
  XNOR2_X1 \Check1_CheckInst_1_U22  ( .A(Red_StateRegOutput[9]), .B(
        Red_SignaltoCheck[137]), .ZN(\Check1_CheckInst_1_n22 ) );
  NOR2_X1 \Check1_CheckInst_1_U21  ( .A1(\Check1_CheckInst_1_n20 ), .A2(
        \Check1_CheckInst_1_n19 ), .ZN(\Check1_CheckInst_1_n28 ) );
  XOR2_X1 \Check1_CheckInst_1_U20  ( .A(Red_Feedback[61]), .B(
        Red_SignaltoCheck[125]), .Z(\Check1_CheckInst_1_n19 ) );
  XOR2_X1 \Check1_CheckInst_1_U19  ( .A(Red_Feedback[53]), .B(
        Red_SignaltoCheck[117]), .Z(\Check1_CheckInst_1_n20 ) );
  NAND2_X1 \Check1_CheckInst_1_U18  ( .A1(\Check1_CheckInst_1_n18 ), .A2(
        \Check1_CheckInst_1_n17 ), .ZN(\Check1_CheckInst_1_n30 ) );
  XNOR2_X1 \Check1_CheckInst_1_U17  ( .A(Red_Feedback[41]), .B(
        Red_SignaltoCheck[105]), .ZN(\Check1_CheckInst_1_n17 ) );
  XNOR2_X1 \Check1_CheckInst_1_U16  ( .A(Red_Feedback[45]), .B(
        Red_SignaltoCheck[109]), .ZN(\Check1_CheckInst_1_n18 ) );
  NAND2_X1 \Check1_CheckInst_1_U15  ( .A1(\Check1_CheckInst_1_n16 ), .A2(
        \Check1_CheckInst_1_n15 ), .ZN(\Check1_CheckInst_1_n96 ) );
  NOR2_X1 \Check1_CheckInst_1_U14  ( .A1(\Check1_CheckInst_1_n14 ), .A2(
        \Check1_CheckInst_1_n13 ), .ZN(\Check1_CheckInst_1_n15 ) );
  NAND2_X1 \Check1_CheckInst_1_U13  ( .A1(\Check1_CheckInst_1_n12 ), .A2(
        \Check1_CheckInst_1_n11 ), .ZN(\Check1_CheckInst_1_n13 ) );
  NOR2_X1 \Check1_CheckInst_1_U12  ( .A1(\Check1_CheckInst_1_n10 ), .A2(
        \Check1_CheckInst_1_n9 ), .ZN(\Check1_CheckInst_1_n11 ) );
  XOR2_X1 \Check1_CheckInst_1_U11  ( .A(Red_Feedback[33]), .B(
        Red_SignaltoCheck[97]), .Z(\Check1_CheckInst_1_n9 ) );
  XOR2_X1 \Check1_CheckInst_1_U10  ( .A(Red_Feedback[49]), .B(
        Red_SignaltoCheck[113]), .Z(\Check1_CheckInst_1_n10 ) );
  NOR2_X1 \Check1_CheckInst_1_U9  ( .A1(\Check1_CheckInst_1_n8 ), .A2(
        \Check1_CheckInst_1_n7 ), .ZN(\Check1_CheckInst_1_n12 ) );
  XOR2_X1 \Check1_CheckInst_1_U8  ( .A(Red_Feedback[37]), .B(
        Red_SignaltoCheck[101]), .Z(\Check1_CheckInst_1_n7 ) );
  XOR2_X1 \Check1_CheckInst_1_U7  ( .A(Red_Feedback[29]), .B(
        Red_SignaltoCheck[93]), .Z(\Check1_CheckInst_1_n8 ) );
  NAND2_X1 \Check1_CheckInst_1_U6  ( .A1(\Check1_CheckInst_1_n6 ), .A2(
        \Check1_CheckInst_1_n5 ), .ZN(\Check1_CheckInst_1_n14 ) );
  XNOR2_X1 \Check1_CheckInst_1_U5  ( .A(Red_StateRegOutput[49]), .B(
        Red_SignaltoCheck[177]), .ZN(\Check1_CheckInst_1_n5 ) );
  XNOR2_X1 \Check1_CheckInst_1_U4  ( .A(Red_StateRegOutput[53]), .B(
        Red_SignaltoCheck[181]), .ZN(\Check1_CheckInst_1_n6 ) );
  NOR2_X1 \Check1_CheckInst_1_U3  ( .A1(\Check1_CheckInst_1_n4 ), .A2(
        \Check1_CheckInst_1_n3 ), .ZN(\Check1_CheckInst_1_n16 ) );
  XOR2_X1 \Check1_CheckInst_1_U2  ( .A(Red_StateRegOutput[41]), .B(
        Red_SignaltoCheck[169]), .Z(\Check1_CheckInst_1_n3 ) );
  XOR2_X1 \Check1_CheckInst_1_U1  ( .A(Red_StateRegOutput[57]), .B(
        Red_SignaltoCheck[185]), .Z(\Check1_CheckInst_1_n4 ) );
  NOR2_X1 \Check1_CheckInst_2_U95  ( .A1(\Check1_CheckInst_2_n96 ), .A2(
        \Check1_CheckInst_2_n95 ), .ZN(Error[2]) );
  NAND2_X1 \Check1_CheckInst_2_U94  ( .A1(\Check1_CheckInst_2_n94 ), .A2(
        \Check1_CheckInst_2_n93 ), .ZN(\Check1_CheckInst_2_n95 ) );
  NOR2_X1 \Check1_CheckInst_2_U93  ( .A1(\Check1_CheckInst_2_n92 ), .A2(
        \Check1_CheckInst_2_n91 ), .ZN(\Check1_CheckInst_2_n93 ) );
  NAND2_X1 \Check1_CheckInst_2_U92  ( .A1(\Check1_CheckInst_2_n90 ), .A2(
        \Check1_CheckInst_2_n89 ), .ZN(\Check1_CheckInst_2_n91 ) );
  NOR2_X1 \Check1_CheckInst_2_U91  ( .A1(\Check1_CheckInst_2_n88 ), .A2(
        \Check1_CheckInst_2_n87 ), .ZN(\Check1_CheckInst_2_n89 ) );
  NAND2_X1 \Check1_CheckInst_2_U90  ( .A1(\Check1_CheckInst_2_n86 ), .A2(
        \Check1_CheckInst_2_n85 ), .ZN(\Check1_CheckInst_2_n87 ) );
  NOR2_X1 \Check1_CheckInst_2_U89  ( .A1(\Check1_CheckInst_2_n84 ), .A2(
        \Check1_CheckInst_2_n83 ), .ZN(\Check1_CheckInst_2_n85 ) );
  NAND2_X1 \Check1_CheckInst_2_U88  ( .A1(\Check1_CheckInst_2_n82 ), .A2(
        \Check1_CheckInst_2_n81 ), .ZN(\Check1_CheckInst_2_n83 ) );
  XNOR2_X1 \Check1_CheckInst_2_U87  ( .A(Red_StateRegOutput[26]), .B(
        Red_SignaltoCheck[154]), .ZN(\Check1_CheckInst_2_n81 ) );
  XNOR2_X1 \Check1_CheckInst_2_U86  ( .A(Red_StateRegOutput[30]), .B(
        Red_SignaltoCheck[158]), .ZN(\Check1_CheckInst_2_n82 ) );
  NAND2_X1 \Check1_CheckInst_2_U85  ( .A1(\Check1_CheckInst_2_n80 ), .A2(
        \Check1_CheckInst_2_n79 ), .ZN(\Check1_CheckInst_2_n84 ) );
  XNOR2_X1 \Check1_CheckInst_2_U84  ( .A(Red_StateRegOutput[46]), .B(
        Red_SignaltoCheck[174]), .ZN(\Check1_CheckInst_2_n79 ) );
  XNOR2_X1 \Check1_CheckInst_2_U83  ( .A(Red_StateRegOutput[38]), .B(
        Red_SignaltoCheck[166]), .ZN(\Check1_CheckInst_2_n80 ) );
  NOR2_X1 \Check1_CheckInst_2_U82  ( .A1(\Check1_CheckInst_2_n78 ), .A2(
        \Check1_CheckInst_2_n77 ), .ZN(\Check1_CheckInst_2_n86 ) );
  NAND2_X1 \Check1_CheckInst_2_U81  ( .A1(\Check1_CheckInst_2_n76 ), .A2(
        \Check1_CheckInst_2_n75 ), .ZN(\Check1_CheckInst_2_n77 ) );
  XNOR2_X1 \Check1_CheckInst_2_U80  ( .A(Red_StateRegOutput[22]), .B(
        Red_SignaltoCheck[150]), .ZN(\Check1_CheckInst_2_n75 ) );
  XNOR2_X1 \Check1_CheckInst_2_U79  ( .A(Red_StateRegOutput[14]), .B(
        Red_SignaltoCheck[142]), .ZN(\Check1_CheckInst_2_n76 ) );
  NAND2_X1 \Check1_CheckInst_2_U78  ( .A1(\Check1_CheckInst_2_n74 ), .A2(
        \Check1_CheckInst_2_n73 ), .ZN(\Check1_CheckInst_2_n78 ) );
  XNOR2_X1 \Check1_CheckInst_2_U77  ( .A(Red_StateRegOutput[18]), .B(
        Red_SignaltoCheck[146]), .ZN(\Check1_CheckInst_2_n73 ) );
  XNOR2_X1 \Check1_CheckInst_2_U76  ( .A(Red_StateRegOutput[34]), .B(
        Red_SignaltoCheck[162]), .ZN(\Check1_CheckInst_2_n74 ) );
  NAND2_X1 \Check1_CheckInst_2_U75  ( .A1(\Check1_CheckInst_2_n72 ), .A2(
        \Check1_CheckInst_2_n71 ), .ZN(\Check1_CheckInst_2_n88 ) );
  NOR2_X1 \Check1_CheckInst_2_U74  ( .A1(\Check1_CheckInst_2_n70 ), .A2(
        \Check1_CheckInst_2_n69 ), .ZN(\Check1_CheckInst_2_n71 ) );
  XOR2_X1 \Check1_CheckInst_2_U73  ( .A(Red_AddRoundKeyOutput[26]), .B(
        Red_SignaltoCheck[26]), .Z(\Check1_CheckInst_2_n69 ) );
  XOR2_X1 \Check1_CheckInst_2_U72  ( .A(Red_AddRoundKeyOutput[42]), .B(
        Red_SignaltoCheck[42]), .Z(\Check1_CheckInst_2_n70 ) );
  NOR2_X1 \Check1_CheckInst_2_U71  ( .A1(\Check1_CheckInst_2_n68 ), .A2(
        \Check1_CheckInst_2_n67 ), .ZN(\Check1_CheckInst_2_n72 ) );
  XOR2_X1 \Check1_CheckInst_2_U70  ( .A(Red_AddRoundKeyOutput[34]), .B(
        Red_SignaltoCheck[34]), .Z(\Check1_CheckInst_2_n67 ) );
  XOR2_X1 \Check1_CheckInst_2_U69  ( .A(Red_AddRoundKeyOutput[38]), .B(
        Red_SignaltoCheck[38]), .Z(\Check1_CheckInst_2_n68 ) );
  NOR2_X1 \Check1_CheckInst_2_U68  ( .A1(\Check1_CheckInst_2_n66 ), .A2(
        \Check1_CheckInst_2_n65 ), .ZN(\Check1_CheckInst_2_n90 ) );
  NAND2_X1 \Check1_CheckInst_2_U67  ( .A1(\Check1_CheckInst_2_n64 ), .A2(
        \Check1_CheckInst_2_n63 ), .ZN(\Check1_CheckInst_2_n65 ) );
  XNOR2_X1 \Check1_CheckInst_2_U66  ( .A(Red_AddRoundKeyOutput[10]), .B(
        Red_SignaltoCheck[10]), .ZN(\Check1_CheckInst_2_n63 ) );
  XNOR2_X1 \Check1_CheckInst_2_U65  ( .A(Red_AddRoundKeyOutput[14]), .B(
        Red_SignaltoCheck[14]), .ZN(\Check1_CheckInst_2_n64 ) );
  NAND2_X1 \Check1_CheckInst_2_U64  ( .A1(\Check1_CheckInst_2_n62 ), .A2(
        \Check1_CheckInst_2_n61 ), .ZN(\Check1_CheckInst_2_n66 ) );
  XNOR2_X1 \Check1_CheckInst_2_U63  ( .A(Red_AddRoundKeyOutput[30]), .B(
        Red_SignaltoCheck[30]), .ZN(\Check1_CheckInst_2_n61 ) );
  XNOR2_X1 \Check1_CheckInst_2_U62  ( .A(Red_AddRoundKeyOutput[22]), .B(
        Red_SignaltoCheck[22]), .ZN(\Check1_CheckInst_2_n62 ) );
  NAND2_X1 \Check1_CheckInst_2_U61  ( .A1(\Check1_CheckInst_2_n60 ), .A2(
        \Check1_CheckInst_2_n59 ), .ZN(\Check1_CheckInst_2_n92 ) );
  NOR2_X1 \Check1_CheckInst_2_U60  ( .A1(\Check1_CheckInst_2_n58 ), .A2(
        \Check1_CheckInst_2_n57 ), .ZN(\Check1_CheckInst_2_n59 ) );
  NAND2_X1 \Check1_CheckInst_2_U59  ( .A1(\Check1_CheckInst_2_n56 ), .A2(
        \Check1_CheckInst_2_n55 ), .ZN(\Check1_CheckInst_2_n57 ) );
  NOR2_X1 \Check1_CheckInst_2_U58  ( .A1(\Check1_CheckInst_2_n54 ), .A2(
        \Check1_CheckInst_2_n53 ), .ZN(\Check1_CheckInst_2_n55 ) );
  NAND2_X1 \Check1_CheckInst_2_U57  ( .A1(\Check1_CheckInst_2_n52 ), .A2(
        \Check1_CheckInst_2_n51 ), .ZN(\Check1_CheckInst_2_n53 ) );
  XNOR2_X1 \Check1_CheckInst_2_U56  ( .A(Red_StateRegOutput[62]), .B(
        Red_SignaltoCheck[190]), .ZN(\Check1_CheckInst_2_n51 ) );
  XNOR2_X1 \Check1_CheckInst_2_U55  ( .A(Red_SignaltoCheck[6]), .B(
        Red_AddRoundKeyOutput[6]), .ZN(\Check1_CheckInst_2_n52 ) );
  NAND2_X1 \Check1_CheckInst_2_U54  ( .A1(\Check1_CheckInst_2_n50 ), .A2(
        \Check1_CheckInst_2_n49 ), .ZN(\Check1_CheckInst_2_n54 ) );
  XNOR2_X1 \Check1_CheckInst_2_U53  ( .A(Red_AddRoundKeyOutput[2]), .B(
        Red_SignaltoCheck[2]), .ZN(\Check1_CheckInst_2_n49 ) );
  XNOR2_X1 \Check1_CheckInst_2_U52  ( .A(Red_AddRoundKeyOutput[18]), .B(
        Red_SignaltoCheck[18]), .ZN(\Check1_CheckInst_2_n50 ) );
  NOR2_X1 \Check1_CheckInst_2_U51  ( .A1(\Check1_CheckInst_2_n48 ), .A2(
        \Check1_CheckInst_2_n47 ), .ZN(\Check1_CheckInst_2_n56 ) );
  NAND2_X1 \Check1_CheckInst_2_U50  ( .A1(\Check1_CheckInst_2_n46 ), .A2(
        \Check1_CheckInst_2_n45 ), .ZN(\Check1_CheckInst_2_n47 ) );
  XNOR2_X1 \Check1_CheckInst_2_U49  ( .A(Red_Feedback[10]), .B(
        Red_SignaltoCheck[74]), .ZN(\Check1_CheckInst_2_n45 ) );
  XNOR2_X1 \Check1_CheckInst_2_U48  ( .A(Red_Feedback[26]), .B(
        Red_SignaltoCheck[90]), .ZN(\Check1_CheckInst_2_n46 ) );
  NAND2_X1 \Check1_CheckInst_2_U47  ( .A1(\Check1_CheckInst_2_n44 ), .A2(
        \Check1_CheckInst_2_n43 ), .ZN(\Check1_CheckInst_2_n48 ) );
  XNOR2_X1 \Check1_CheckInst_2_U46  ( .A(Red_Feedback[18]), .B(
        Red_SignaltoCheck[82]), .ZN(\Check1_CheckInst_2_n43 ) );
  XNOR2_X1 \Check1_CheckInst_2_U45  ( .A(Red_Feedback[22]), .B(
        Red_SignaltoCheck[86]), .ZN(\Check1_CheckInst_2_n44 ) );
  NAND2_X1 \Check1_CheckInst_2_U44  ( .A1(\Check1_CheckInst_2_n42 ), .A2(
        \Check1_CheckInst_2_n41 ), .ZN(\Check1_CheckInst_2_n58 ) );
  NOR2_X1 \Check1_CheckInst_2_U43  ( .A1(\Check1_CheckInst_2_n40 ), .A2(
        \Check1_CheckInst_2_n39 ), .ZN(\Check1_CheckInst_2_n41 ) );
  XOR2_X1 \Check1_CheckInst_2_U42  ( .A(Red_AddRoundKeyOutput[58]), .B(
        Red_SignaltoCheck[58]), .Z(\Check1_CheckInst_2_n39 ) );
  XOR2_X1 \Check1_CheckInst_2_U41  ( .A(Red_AddRoundKeyOutput[62]), .B(
        Red_SignaltoCheck[62]), .Z(\Check1_CheckInst_2_n40 ) );
  NOR2_X1 \Check1_CheckInst_2_U40  ( .A1(\Check1_CheckInst_2_n38 ), .A2(
        \Check1_CheckInst_2_n37 ), .ZN(\Check1_CheckInst_2_n42 ) );
  XOR2_X1 \Check1_CheckInst_2_U39  ( .A(Red_Feedback[14]), .B(
        Red_SignaltoCheck[78]), .Z(\Check1_CheckInst_2_n37 ) );
  XOR2_X1 \Check1_CheckInst_2_U38  ( .A(Red_Feedback[6]), .B(
        Red_SignaltoCheck[70]), .Z(\Check1_CheckInst_2_n38 ) );
  NOR2_X1 \Check1_CheckInst_2_U37  ( .A1(\Check1_CheckInst_2_n36 ), .A2(
        \Check1_CheckInst_2_n35 ), .ZN(\Check1_CheckInst_2_n60 ) );
  NAND2_X1 \Check1_CheckInst_2_U36  ( .A1(\Check1_CheckInst_2_n34 ), .A2(
        \Check1_CheckInst_2_n33 ), .ZN(\Check1_CheckInst_2_n35 ) );
  XNOR2_X1 \Check1_CheckInst_2_U35  ( .A(Red_AddRoundKeyOutput[54]), .B(
        Red_SignaltoCheck[54]), .ZN(\Check1_CheckInst_2_n33 ) );
  XNOR2_X1 \Check1_CheckInst_2_U34  ( .A(Red_AddRoundKeyOutput[46]), .B(
        Red_SignaltoCheck[46]), .ZN(\Check1_CheckInst_2_n34 ) );
  NAND2_X1 \Check1_CheckInst_2_U33  ( .A1(\Check1_CheckInst_2_n32 ), .A2(
        \Check1_CheckInst_2_n31 ), .ZN(\Check1_CheckInst_2_n36 ) );
  XNOR2_X1 \Check1_CheckInst_2_U32  ( .A(Red_AddRoundKeyOutput[50]), .B(
        Red_SignaltoCheck[50]), .ZN(\Check1_CheckInst_2_n31 ) );
  XNOR2_X1 \Check1_CheckInst_2_U31  ( .A(Red_Feedback[2]), .B(
        Red_SignaltoCheck[66]), .ZN(\Check1_CheckInst_2_n32 ) );
  NOR2_X1 \Check1_CheckInst_2_U30  ( .A1(\Check1_CheckInst_2_n30 ), .A2(
        \Check1_CheckInst_2_n29 ), .ZN(\Check1_CheckInst_2_n94 ) );
  NAND2_X1 \Check1_CheckInst_2_U29  ( .A1(\Check1_CheckInst_2_n28 ), .A2(
        \Check1_CheckInst_2_n27 ), .ZN(\Check1_CheckInst_2_n29 ) );
  NOR2_X1 \Check1_CheckInst_2_U28  ( .A1(\Check1_CheckInst_2_n26 ), .A2(
        \Check1_CheckInst_2_n25 ), .ZN(\Check1_CheckInst_2_n27 ) );
  NAND2_X1 \Check1_CheckInst_2_U27  ( .A1(\Check1_CheckInst_2_n24 ), .A2(
        \Check1_CheckInst_2_n23 ), .ZN(\Check1_CheckInst_2_n25 ) );
  XNOR2_X1 \Check1_CheckInst_2_U26  ( .A(Red_StateRegOutput[2]), .B(
        Red_SignaltoCheck[130]), .ZN(\Check1_CheckInst_2_n23 ) );
  XNOR2_X1 \Check1_CheckInst_2_U25  ( .A(Red_StateRegOutput[6]), .B(
        Red_SignaltoCheck[134]), .ZN(\Check1_CheckInst_2_n24 ) );
  NAND2_X1 \Check1_CheckInst_2_U24  ( .A1(\Check1_CheckInst_2_n22 ), .A2(
        \Check1_CheckInst_2_n21 ), .ZN(\Check1_CheckInst_2_n26 ) );
  XNOR2_X1 \Check1_CheckInst_2_U23  ( .A(Red_Feedback[58]), .B(
        Red_SignaltoCheck[122]), .ZN(\Check1_CheckInst_2_n21 ) );
  XNOR2_X1 \Check1_CheckInst_2_U22  ( .A(Red_StateRegOutput[10]), .B(
        Red_SignaltoCheck[138]), .ZN(\Check1_CheckInst_2_n22 ) );
  NOR2_X1 \Check1_CheckInst_2_U21  ( .A1(\Check1_CheckInst_2_n20 ), .A2(
        \Check1_CheckInst_2_n19 ), .ZN(\Check1_CheckInst_2_n28 ) );
  XOR2_X1 \Check1_CheckInst_2_U20  ( .A(Red_Feedback[62]), .B(
        Red_SignaltoCheck[126]), .Z(\Check1_CheckInst_2_n19 ) );
  XOR2_X1 \Check1_CheckInst_2_U19  ( .A(Red_Feedback[54]), .B(
        Red_SignaltoCheck[118]), .Z(\Check1_CheckInst_2_n20 ) );
  NAND2_X1 \Check1_CheckInst_2_U18  ( .A1(\Check1_CheckInst_2_n18 ), .A2(
        \Check1_CheckInst_2_n17 ), .ZN(\Check1_CheckInst_2_n30 ) );
  XNOR2_X1 \Check1_CheckInst_2_U17  ( .A(Red_Feedback[42]), .B(
        Red_SignaltoCheck[106]), .ZN(\Check1_CheckInst_2_n17 ) );
  XNOR2_X1 \Check1_CheckInst_2_U16  ( .A(Red_Feedback[46]), .B(
        Red_SignaltoCheck[110]), .ZN(\Check1_CheckInst_2_n18 ) );
  NAND2_X1 \Check1_CheckInst_2_U15  ( .A1(\Check1_CheckInst_2_n16 ), .A2(
        \Check1_CheckInst_2_n15 ), .ZN(\Check1_CheckInst_2_n96 ) );
  NOR2_X1 \Check1_CheckInst_2_U14  ( .A1(\Check1_CheckInst_2_n14 ), .A2(
        \Check1_CheckInst_2_n13 ), .ZN(\Check1_CheckInst_2_n15 ) );
  NAND2_X1 \Check1_CheckInst_2_U13  ( .A1(\Check1_CheckInst_2_n12 ), .A2(
        \Check1_CheckInst_2_n11 ), .ZN(\Check1_CheckInst_2_n13 ) );
  NOR2_X1 \Check1_CheckInst_2_U12  ( .A1(\Check1_CheckInst_2_n10 ), .A2(
        \Check1_CheckInst_2_n9 ), .ZN(\Check1_CheckInst_2_n11 ) );
  XOR2_X1 \Check1_CheckInst_2_U11  ( .A(Red_Feedback[34]), .B(
        Red_SignaltoCheck[98]), .Z(\Check1_CheckInst_2_n9 ) );
  XOR2_X1 \Check1_CheckInst_2_U10  ( .A(Red_Feedback[50]), .B(
        Red_SignaltoCheck[114]), .Z(\Check1_CheckInst_2_n10 ) );
  NOR2_X1 \Check1_CheckInst_2_U9  ( .A1(\Check1_CheckInst_2_n8 ), .A2(
        \Check1_CheckInst_2_n7 ), .ZN(\Check1_CheckInst_2_n12 ) );
  XOR2_X1 \Check1_CheckInst_2_U8  ( .A(Red_Feedback[38]), .B(
        Red_SignaltoCheck[102]), .Z(\Check1_CheckInst_2_n7 ) );
  XOR2_X1 \Check1_CheckInst_2_U7  ( .A(Red_Feedback[30]), .B(
        Red_SignaltoCheck[94]), .Z(\Check1_CheckInst_2_n8 ) );
  NAND2_X1 \Check1_CheckInst_2_U6  ( .A1(\Check1_CheckInst_2_n6 ), .A2(
        \Check1_CheckInst_2_n5 ), .ZN(\Check1_CheckInst_2_n14 ) );
  XNOR2_X1 \Check1_CheckInst_2_U5  ( .A(Red_StateRegOutput[50]), .B(
        Red_SignaltoCheck[178]), .ZN(\Check1_CheckInst_2_n5 ) );
  XNOR2_X1 \Check1_CheckInst_2_U4  ( .A(Red_StateRegOutput[54]), .B(
        Red_SignaltoCheck[182]), .ZN(\Check1_CheckInst_2_n6 ) );
  NOR2_X1 \Check1_CheckInst_2_U3  ( .A1(\Check1_CheckInst_2_n4 ), .A2(
        \Check1_CheckInst_2_n3 ), .ZN(\Check1_CheckInst_2_n16 ) );
  XOR2_X1 \Check1_CheckInst_2_U2  ( .A(Red_StateRegOutput[42]), .B(
        Red_SignaltoCheck[170]), .Z(\Check1_CheckInst_2_n3 ) );
  XOR2_X1 \Check1_CheckInst_2_U1  ( .A(Red_StateRegOutput[58]), .B(
        Red_SignaltoCheck[186]), .Z(\Check1_CheckInst_2_n4 ) );
  NOR2_X1 \Check1_CheckInst_3_U95  ( .A1(\Check1_CheckInst_3_n96 ), .A2(
        \Check1_CheckInst_3_n95 ), .ZN(Error[3]) );
  NAND2_X1 \Check1_CheckInst_3_U94  ( .A1(\Check1_CheckInst_3_n94 ), .A2(
        \Check1_CheckInst_3_n93 ), .ZN(\Check1_CheckInst_3_n95 ) );
  NOR2_X1 \Check1_CheckInst_3_U93  ( .A1(\Check1_CheckInst_3_n92 ), .A2(
        \Check1_CheckInst_3_n91 ), .ZN(\Check1_CheckInst_3_n93 ) );
  NAND2_X1 \Check1_CheckInst_3_U92  ( .A1(\Check1_CheckInst_3_n90 ), .A2(
        \Check1_CheckInst_3_n89 ), .ZN(\Check1_CheckInst_3_n91 ) );
  NOR2_X1 \Check1_CheckInst_3_U91  ( .A1(\Check1_CheckInst_3_n88 ), .A2(
        \Check1_CheckInst_3_n87 ), .ZN(\Check1_CheckInst_3_n89 ) );
  NAND2_X1 \Check1_CheckInst_3_U90  ( .A1(\Check1_CheckInst_3_n86 ), .A2(
        \Check1_CheckInst_3_n85 ), .ZN(\Check1_CheckInst_3_n87 ) );
  NOR2_X1 \Check1_CheckInst_3_U89  ( .A1(\Check1_CheckInst_3_n84 ), .A2(
        \Check1_CheckInst_3_n83 ), .ZN(\Check1_CheckInst_3_n85 ) );
  NAND2_X1 \Check1_CheckInst_3_U88  ( .A1(\Check1_CheckInst_3_n82 ), .A2(
        \Check1_CheckInst_3_n81 ), .ZN(\Check1_CheckInst_3_n83 ) );
  XNOR2_X1 \Check1_CheckInst_3_U87  ( .A(Red_StateRegOutput[27]), .B(
        Red_SignaltoCheck[155]), .ZN(\Check1_CheckInst_3_n81 ) );
  XNOR2_X1 \Check1_CheckInst_3_U86  ( .A(Red_StateRegOutput[31]), .B(
        Red_SignaltoCheck[159]), .ZN(\Check1_CheckInst_3_n82 ) );
  NAND2_X1 \Check1_CheckInst_3_U85  ( .A1(\Check1_CheckInst_3_n80 ), .A2(
        \Check1_CheckInst_3_n79 ), .ZN(\Check1_CheckInst_3_n84 ) );
  XNOR2_X1 \Check1_CheckInst_3_U84  ( .A(Red_StateRegOutput[47]), .B(
        Red_SignaltoCheck[175]), .ZN(\Check1_CheckInst_3_n79 ) );
  XNOR2_X1 \Check1_CheckInst_3_U83  ( .A(Red_StateRegOutput[39]), .B(
        Red_SignaltoCheck[167]), .ZN(\Check1_CheckInst_3_n80 ) );
  NOR2_X1 \Check1_CheckInst_3_U82  ( .A1(\Check1_CheckInst_3_n78 ), .A2(
        \Check1_CheckInst_3_n77 ), .ZN(\Check1_CheckInst_3_n86 ) );
  NAND2_X1 \Check1_CheckInst_3_U81  ( .A1(\Check1_CheckInst_3_n76 ), .A2(
        \Check1_CheckInst_3_n75 ), .ZN(\Check1_CheckInst_3_n77 ) );
  XNOR2_X1 \Check1_CheckInst_3_U80  ( .A(Red_StateRegOutput[23]), .B(
        Red_SignaltoCheck[151]), .ZN(\Check1_CheckInst_3_n75 ) );
  XNOR2_X1 \Check1_CheckInst_3_U79  ( .A(Red_StateRegOutput[15]), .B(
        Red_SignaltoCheck[143]), .ZN(\Check1_CheckInst_3_n76 ) );
  NAND2_X1 \Check1_CheckInst_3_U78  ( .A1(\Check1_CheckInst_3_n74 ), .A2(
        \Check1_CheckInst_3_n73 ), .ZN(\Check1_CheckInst_3_n78 ) );
  XNOR2_X1 \Check1_CheckInst_3_U77  ( .A(Red_StateRegOutput[19]), .B(
        Red_SignaltoCheck[147]), .ZN(\Check1_CheckInst_3_n73 ) );
  XNOR2_X1 \Check1_CheckInst_3_U76  ( .A(Red_StateRegOutput[35]), .B(
        Red_SignaltoCheck[163]), .ZN(\Check1_CheckInst_3_n74 ) );
  NAND2_X1 \Check1_CheckInst_3_U75  ( .A1(\Check1_CheckInst_3_n72 ), .A2(
        \Check1_CheckInst_3_n71 ), .ZN(\Check1_CheckInst_3_n88 ) );
  NOR2_X1 \Check1_CheckInst_3_U74  ( .A1(\Check1_CheckInst_3_n70 ), .A2(
        \Check1_CheckInst_3_n69 ), .ZN(\Check1_CheckInst_3_n71 ) );
  XOR2_X1 \Check1_CheckInst_3_U73  ( .A(Red_AddRoundKeyOutput[27]), .B(
        Red_SignaltoCheck[27]), .Z(\Check1_CheckInst_3_n69 ) );
  XOR2_X1 \Check1_CheckInst_3_U72  ( .A(Red_AddRoundKeyOutput[43]), .B(
        Red_SignaltoCheck[43]), .Z(\Check1_CheckInst_3_n70 ) );
  NOR2_X1 \Check1_CheckInst_3_U71  ( .A1(\Check1_CheckInst_3_n68 ), .A2(
        \Check1_CheckInst_3_n67 ), .ZN(\Check1_CheckInst_3_n72 ) );
  XOR2_X1 \Check1_CheckInst_3_U70  ( .A(Red_AddRoundKeyOutput[35]), .B(
        Red_SignaltoCheck[35]), .Z(\Check1_CheckInst_3_n67 ) );
  XOR2_X1 \Check1_CheckInst_3_U69  ( .A(Red_AddRoundKeyOutput[39]), .B(
        Red_SignaltoCheck[39]), .Z(\Check1_CheckInst_3_n68 ) );
  NOR2_X1 \Check1_CheckInst_3_U68  ( .A1(\Check1_CheckInst_3_n66 ), .A2(
        \Check1_CheckInst_3_n65 ), .ZN(\Check1_CheckInst_3_n90 ) );
  NAND2_X1 \Check1_CheckInst_3_U67  ( .A1(\Check1_CheckInst_3_n64 ), .A2(
        \Check1_CheckInst_3_n63 ), .ZN(\Check1_CheckInst_3_n65 ) );
  XNOR2_X1 \Check1_CheckInst_3_U66  ( .A(Red_AddRoundKeyOutput[11]), .B(
        Red_SignaltoCheck[11]), .ZN(\Check1_CheckInst_3_n63 ) );
  XNOR2_X1 \Check1_CheckInst_3_U65  ( .A(Red_AddRoundKeyOutput[15]), .B(
        Red_SignaltoCheck[15]), .ZN(\Check1_CheckInst_3_n64 ) );
  NAND2_X1 \Check1_CheckInst_3_U64  ( .A1(\Check1_CheckInst_3_n62 ), .A2(
        \Check1_CheckInst_3_n61 ), .ZN(\Check1_CheckInst_3_n66 ) );
  XNOR2_X1 \Check1_CheckInst_3_U63  ( .A(Red_AddRoundKeyOutput[31]), .B(
        Red_SignaltoCheck[31]), .ZN(\Check1_CheckInst_3_n61 ) );
  XNOR2_X1 \Check1_CheckInst_3_U62  ( .A(Red_AddRoundKeyOutput[23]), .B(
        Red_SignaltoCheck[23]), .ZN(\Check1_CheckInst_3_n62 ) );
  NAND2_X1 \Check1_CheckInst_3_U61  ( .A1(\Check1_CheckInst_3_n60 ), .A2(
        \Check1_CheckInst_3_n59 ), .ZN(\Check1_CheckInst_3_n92 ) );
  NOR2_X1 \Check1_CheckInst_3_U60  ( .A1(\Check1_CheckInst_3_n58 ), .A2(
        \Check1_CheckInst_3_n57 ), .ZN(\Check1_CheckInst_3_n59 ) );
  NAND2_X1 \Check1_CheckInst_3_U59  ( .A1(\Check1_CheckInst_3_n56 ), .A2(
        \Check1_CheckInst_3_n55 ), .ZN(\Check1_CheckInst_3_n57 ) );
  NOR2_X1 \Check1_CheckInst_3_U58  ( .A1(\Check1_CheckInst_3_n54 ), .A2(
        \Check1_CheckInst_3_n53 ), .ZN(\Check1_CheckInst_3_n55 ) );
  NAND2_X1 \Check1_CheckInst_3_U57  ( .A1(\Check1_CheckInst_3_n52 ), .A2(
        \Check1_CheckInst_3_n51 ), .ZN(\Check1_CheckInst_3_n53 ) );
  XNOR2_X1 \Check1_CheckInst_3_U56  ( .A(Red_StateRegOutput[63]), .B(
        Red_SignaltoCheck[191]), .ZN(\Check1_CheckInst_3_n51 ) );
  XNOR2_X1 \Check1_CheckInst_3_U55  ( .A(Red_SignaltoCheck[7]), .B(
        Red_AddRoundKeyOutput[7]), .ZN(\Check1_CheckInst_3_n52 ) );
  NAND2_X1 \Check1_CheckInst_3_U54  ( .A1(\Check1_CheckInst_3_n50 ), .A2(
        \Check1_CheckInst_3_n49 ), .ZN(\Check1_CheckInst_3_n54 ) );
  XNOR2_X1 \Check1_CheckInst_3_U53  ( .A(Red_AddRoundKeyOutput[3]), .B(
        Red_SignaltoCheck[3]), .ZN(\Check1_CheckInst_3_n49 ) );
  XNOR2_X1 \Check1_CheckInst_3_U52  ( .A(Red_AddRoundKeyOutput[19]), .B(
        Red_SignaltoCheck[19]), .ZN(\Check1_CheckInst_3_n50 ) );
  NOR2_X1 \Check1_CheckInst_3_U51  ( .A1(\Check1_CheckInst_3_n48 ), .A2(
        \Check1_CheckInst_3_n47 ), .ZN(\Check1_CheckInst_3_n56 ) );
  NAND2_X1 \Check1_CheckInst_3_U50  ( .A1(\Check1_CheckInst_3_n46 ), .A2(
        \Check1_CheckInst_3_n45 ), .ZN(\Check1_CheckInst_3_n47 ) );
  XNOR2_X1 \Check1_CheckInst_3_U49  ( .A(Red_Feedback[11]), .B(
        Red_SignaltoCheck[75]), .ZN(\Check1_CheckInst_3_n45 ) );
  XNOR2_X1 \Check1_CheckInst_3_U48  ( .A(Red_Feedback[27]), .B(
        Red_SignaltoCheck[91]), .ZN(\Check1_CheckInst_3_n46 ) );
  NAND2_X1 \Check1_CheckInst_3_U47  ( .A1(\Check1_CheckInst_3_n44 ), .A2(
        \Check1_CheckInst_3_n43 ), .ZN(\Check1_CheckInst_3_n48 ) );
  XNOR2_X1 \Check1_CheckInst_3_U46  ( .A(Red_Feedback[19]), .B(
        Red_SignaltoCheck[83]), .ZN(\Check1_CheckInst_3_n43 ) );
  XNOR2_X1 \Check1_CheckInst_3_U45  ( .A(Red_Feedback[23]), .B(
        Red_SignaltoCheck[87]), .ZN(\Check1_CheckInst_3_n44 ) );
  NAND2_X1 \Check1_CheckInst_3_U44  ( .A1(\Check1_CheckInst_3_n42 ), .A2(
        \Check1_CheckInst_3_n41 ), .ZN(\Check1_CheckInst_3_n58 ) );
  NOR2_X1 \Check1_CheckInst_3_U43  ( .A1(\Check1_CheckInst_3_n40 ), .A2(
        \Check1_CheckInst_3_n39 ), .ZN(\Check1_CheckInst_3_n41 ) );
  XOR2_X1 \Check1_CheckInst_3_U42  ( .A(Red_AddRoundKeyOutput[59]), .B(
        Red_SignaltoCheck[59]), .Z(\Check1_CheckInst_3_n39 ) );
  XOR2_X1 \Check1_CheckInst_3_U41  ( .A(Red_AddRoundKeyOutput[63]), .B(
        Red_SignaltoCheck[63]), .Z(\Check1_CheckInst_3_n40 ) );
  NOR2_X1 \Check1_CheckInst_3_U40  ( .A1(\Check1_CheckInst_3_n38 ), .A2(
        \Check1_CheckInst_3_n37 ), .ZN(\Check1_CheckInst_3_n42 ) );
  XOR2_X1 \Check1_CheckInst_3_U39  ( .A(Red_Feedback[15]), .B(
        Red_SignaltoCheck[79]), .Z(\Check1_CheckInst_3_n37 ) );
  XOR2_X1 \Check1_CheckInst_3_U38  ( .A(Red_Feedback[7]), .B(
        Red_SignaltoCheck[71]), .Z(\Check1_CheckInst_3_n38 ) );
  NOR2_X1 \Check1_CheckInst_3_U37  ( .A1(\Check1_CheckInst_3_n36 ), .A2(
        \Check1_CheckInst_3_n35 ), .ZN(\Check1_CheckInst_3_n60 ) );
  NAND2_X1 \Check1_CheckInst_3_U36  ( .A1(\Check1_CheckInst_3_n34 ), .A2(
        \Check1_CheckInst_3_n33 ), .ZN(\Check1_CheckInst_3_n35 ) );
  XNOR2_X1 \Check1_CheckInst_3_U35  ( .A(Red_AddRoundKeyOutput[55]), .B(
        Red_SignaltoCheck[55]), .ZN(\Check1_CheckInst_3_n33 ) );
  XNOR2_X1 \Check1_CheckInst_3_U34  ( .A(Red_AddRoundKeyOutput[47]), .B(
        Red_SignaltoCheck[47]), .ZN(\Check1_CheckInst_3_n34 ) );
  NAND2_X1 \Check1_CheckInst_3_U33  ( .A1(\Check1_CheckInst_3_n32 ), .A2(
        \Check1_CheckInst_3_n31 ), .ZN(\Check1_CheckInst_3_n36 ) );
  XNOR2_X1 \Check1_CheckInst_3_U32  ( .A(Red_AddRoundKeyOutput[51]), .B(
        Red_SignaltoCheck[51]), .ZN(\Check1_CheckInst_3_n31 ) );
  XNOR2_X1 \Check1_CheckInst_3_U31  ( .A(Red_Feedback[3]), .B(
        Red_SignaltoCheck[67]), .ZN(\Check1_CheckInst_3_n32 ) );
  NOR2_X1 \Check1_CheckInst_3_U30  ( .A1(\Check1_CheckInst_3_n30 ), .A2(
        \Check1_CheckInst_3_n29 ), .ZN(\Check1_CheckInst_3_n94 ) );
  NAND2_X1 \Check1_CheckInst_3_U29  ( .A1(\Check1_CheckInst_3_n28 ), .A2(
        \Check1_CheckInst_3_n27 ), .ZN(\Check1_CheckInst_3_n29 ) );
  NOR2_X1 \Check1_CheckInst_3_U28  ( .A1(\Check1_CheckInst_3_n26 ), .A2(
        \Check1_CheckInst_3_n25 ), .ZN(\Check1_CheckInst_3_n27 ) );
  NAND2_X1 \Check1_CheckInst_3_U27  ( .A1(\Check1_CheckInst_3_n24 ), .A2(
        \Check1_CheckInst_3_n23 ), .ZN(\Check1_CheckInst_3_n25 ) );
  XNOR2_X1 \Check1_CheckInst_3_U26  ( .A(Red_StateRegOutput[3]), .B(
        Red_SignaltoCheck[131]), .ZN(\Check1_CheckInst_3_n23 ) );
  XNOR2_X1 \Check1_CheckInst_3_U25  ( .A(Red_StateRegOutput[7]), .B(
        Red_SignaltoCheck[135]), .ZN(\Check1_CheckInst_3_n24 ) );
  NAND2_X1 \Check1_CheckInst_3_U24  ( .A1(\Check1_CheckInst_3_n22 ), .A2(
        \Check1_CheckInst_3_n21 ), .ZN(\Check1_CheckInst_3_n26 ) );
  XNOR2_X1 \Check1_CheckInst_3_U23  ( .A(Red_Feedback[59]), .B(
        Red_SignaltoCheck[123]), .ZN(\Check1_CheckInst_3_n21 ) );
  XNOR2_X1 \Check1_CheckInst_3_U22  ( .A(Red_StateRegOutput[11]), .B(
        Red_SignaltoCheck[139]), .ZN(\Check1_CheckInst_3_n22 ) );
  NOR2_X1 \Check1_CheckInst_3_U21  ( .A1(\Check1_CheckInst_3_n20 ), .A2(
        \Check1_CheckInst_3_n19 ), .ZN(\Check1_CheckInst_3_n28 ) );
  XOR2_X1 \Check1_CheckInst_3_U20  ( .A(Red_Feedback[63]), .B(
        Red_SignaltoCheck[127]), .Z(\Check1_CheckInst_3_n19 ) );
  XOR2_X1 \Check1_CheckInst_3_U19  ( .A(Red_Feedback[55]), .B(
        Red_SignaltoCheck[119]), .Z(\Check1_CheckInst_3_n20 ) );
  NAND2_X1 \Check1_CheckInst_3_U18  ( .A1(\Check1_CheckInst_3_n18 ), .A2(
        \Check1_CheckInst_3_n17 ), .ZN(\Check1_CheckInst_3_n30 ) );
  XNOR2_X1 \Check1_CheckInst_3_U17  ( .A(Red_Feedback[43]), .B(
        Red_SignaltoCheck[107]), .ZN(\Check1_CheckInst_3_n17 ) );
  XNOR2_X1 \Check1_CheckInst_3_U16  ( .A(Red_Feedback[47]), .B(
        Red_SignaltoCheck[111]), .ZN(\Check1_CheckInst_3_n18 ) );
  NAND2_X1 \Check1_CheckInst_3_U15  ( .A1(\Check1_CheckInst_3_n16 ), .A2(
        \Check1_CheckInst_3_n15 ), .ZN(\Check1_CheckInst_3_n96 ) );
  NOR2_X1 \Check1_CheckInst_3_U14  ( .A1(\Check1_CheckInst_3_n14 ), .A2(
        \Check1_CheckInst_3_n13 ), .ZN(\Check1_CheckInst_3_n15 ) );
  NAND2_X1 \Check1_CheckInst_3_U13  ( .A1(\Check1_CheckInst_3_n12 ), .A2(
        \Check1_CheckInst_3_n11 ), .ZN(\Check1_CheckInst_3_n13 ) );
  NOR2_X1 \Check1_CheckInst_3_U12  ( .A1(\Check1_CheckInst_3_n10 ), .A2(
        \Check1_CheckInst_3_n9 ), .ZN(\Check1_CheckInst_3_n11 ) );
  XOR2_X1 \Check1_CheckInst_3_U11  ( .A(Red_Feedback[35]), .B(
        Red_SignaltoCheck[99]), .Z(\Check1_CheckInst_3_n9 ) );
  XOR2_X1 \Check1_CheckInst_3_U10  ( .A(Red_Feedback[51]), .B(
        Red_SignaltoCheck[115]), .Z(\Check1_CheckInst_3_n10 ) );
  NOR2_X1 \Check1_CheckInst_3_U9  ( .A1(\Check1_CheckInst_3_n8 ), .A2(
        \Check1_CheckInst_3_n7 ), .ZN(\Check1_CheckInst_3_n12 ) );
  XOR2_X1 \Check1_CheckInst_3_U8  ( .A(Red_Feedback[39]), .B(
        Red_SignaltoCheck[103]), .Z(\Check1_CheckInst_3_n7 ) );
  XOR2_X1 \Check1_CheckInst_3_U7  ( .A(Red_Feedback[31]), .B(
        Red_SignaltoCheck[95]), .Z(\Check1_CheckInst_3_n8 ) );
  NAND2_X1 \Check1_CheckInst_3_U6  ( .A1(\Check1_CheckInst_3_n6 ), .A2(
        \Check1_CheckInst_3_n5 ), .ZN(\Check1_CheckInst_3_n14 ) );
  XNOR2_X1 \Check1_CheckInst_3_U5  ( .A(Red_StateRegOutput[51]), .B(
        Red_SignaltoCheck[179]), .ZN(\Check1_CheckInst_3_n5 ) );
  XNOR2_X1 \Check1_CheckInst_3_U4  ( .A(Red_StateRegOutput[55]), .B(
        Red_SignaltoCheck[183]), .ZN(\Check1_CheckInst_3_n6 ) );
  NOR2_X1 \Check1_CheckInst_3_U3  ( .A1(\Check1_CheckInst_3_n4 ), .A2(
        \Check1_CheckInst_3_n3 ), .ZN(\Check1_CheckInst_3_n16 ) );
  XOR2_X1 \Check1_CheckInst_3_U2  ( .A(Red_StateRegOutput[43]), .B(
        Red_SignaltoCheck[171]), .Z(\Check1_CheckInst_3_n3 ) );
  XOR2_X1 \Check1_CheckInst_3_U1  ( .A(Red_StateRegOutput[59]), .B(
        Red_SignaltoCheck[187]), .Z(\Check1_CheckInst_3_n4 ) );
endmodule

